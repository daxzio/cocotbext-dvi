//
//Written by GowinSynthesis
//Product Version "GowinSynthesis V1.9.7.02Beta"
//Thu Feb 25 16:22:41 2021

//Source file index table:
//file0 "\D:/Gowin/Gowin_V1.9.7.02Beta/IDE/ipcore/DVI_TX/data/dvi_tx_top.v"
//file1 "\D:/Gowin/Gowin_V1.9.7.02Beta/IDE/ipcore/DVI_TX/data/rgb2dvi.vp"
`timescale 100 ps/100 ps
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity",key_keyname="SYNP05_001",key_method="rsa"
`pragma protect key_block
U0dw3aYFMouH3CXEDfA6e/cdu9VXSxccK8hIIFERzi82ZqxoGn6nQL4D6R4O5q/+CErnyvQPKgb2
dATLwZUhnrhlzTJKbmvMljyK7GiaENbwstS1oql6oPHIQvCUyX6Ou3XRaG7ZGOfVRqNPvSrd8Yod
J5MOPRb7naSIietIk29pdfkDofyf7KK8Y1impOPHLYK2ug5Os3N++K4nifldA0kKXJfrGIO5tUwK
uaYKm3pHrKUGR72R2cAfEYSg9EJSSXKziyG+VVoYfagzj5tyqDQPlA9eXw24FUXZBu5qPN5C5i/C
xzrBIahP5ha0mqcHu37qwFuePWJNGYM8NgN9Ig==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin",key_keyname="GoWin001",key_method="rsa"
`pragma protect key_block
coQEjeeFBiYzfVU89oj5lF110E4FutGS+KE/zevm0VJsKRFp99UHVUK56DD7mJegkO/CZ/0xMfYX
OwtzYkiExdGVwHjtyucZpz7HyhyDrJIeLxhUZzo/6RN3axIztxHCmAab64CWC+tUrrgZ6UZZsYEJ
SqrRSJRLtikxqvRYv62hd+UApsl6YyY/NdUmhFrWzh+cA1xO3xKsITEcAg5E/cqiDmkP1BH3/0+F
m4TtYiiu4UxZDQdzz8Ey10T1hP9Y9qvl8uQD2baJF7aVFHTUFaRrqaz/XN+uuL6rm7TJcyoMzAEN
QazMw/gxVQN8++Q+nNsr4Oi9Ka3JtISK77fncw==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=59296)
`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
fC7HWzXWlOj3lIyq7jVYeY5PFx5QpdjytqRjX2ljkIqQwCADPnl0+ilx14F1AoSX3/l3qAWET5Vs
K3ErGGAd2Q3EMfKrb/G7PsdkixiBHoiU5sEkCQYuG5DbTzA9Xs9zsqr8AtEgHujydag1++m5cT9+
Odk86keVwn+oecJlMAS6OP3n/SDWpieX7gQ8jwuciXPvIpQJjdRf/w/9uVaMdai99YEh0jjLHpPT
hM5cNghxHleLKbdS3rXzG0Io8ddpuO8uaJ9E8RVTzcbAs0RVyElC3+FiuClOWEns+KE4KzK72Fql
eDdTIYvmIJ1WXtKJGBsCvS0QSTtQcnHama6wRUt28WE4NBkVrF1RIpV0ZGfqA7paQ0S5tQSXcmgw
K7FN0WsCdKPq9jqds9eL72ZNNhG2v4+YF/NLIzLTrka7uDK8dg84pMGZG+sEeaMzoq2rtAkN0JyE
JuGB0uzNYc+E1XlNQxSVIvKzTT6YTEbcR/6sER0oex8NjHuWodqhb0ufDm9D3/2ow8XZyxgpxOnv
1ye6k1KJDf2L09kiLgGW9HvZAYjhLb1QmNWRKFFnHiXa2yGnodlR/PAcoP6GG+RYG8qYe9BR82Tg
/HIvRRVa6KkKztna2C5dMCBp98SvecOp9BZxu6mSv5b/+gAKq/DQaWf+7XFCsEZrF/b5mIAI9dWL
+ZUGnG0elre3MHcgBljs+a6xNsdv/MTA7EIs4y4yHzgbICDjgKFGOGVSO/tl8JJnRAy1dilDKsKR
tuzew0zOYeheaE5W7cmOuKBhhcD5OaNyF7+eLC40ePx/fqT6mGD8W7J9zhCj4ZPxFzkQzuw+TFdz
2dU4cuzg1nOCZghZ4V64UQXa6bpE4decAy+Ks+tIYwaLhvMmmPLiGURYJB1nUXV9TtCk9bul/GL9
rC1klWdFkJJncXhyBx+ZhVs7uwq+zaUr4eFpCTueo74S8u/F2BrtHHRh64/3P534NIyxVbdfsu9C
EGy7ScwxxrQ5q+TRWBBAQqwpQqQuocsPml8LmL02BvmHctAj0f5wPobXVx53I57BBOdQOMM21W8I
gcFvgoLYWvwvheFBu7pAtaDPpo1QUYpc+fY/7spbWqnHqfC3++9gKCBszQ5pbLmYHRowPs+ujP/d
Z8K/tU9363wez3OL7IuMHGgV7vasWE+KbH8TSRStpKnWlKa0d6TyuAjqcfOGKM2W6jjcno5+4OfH
6fmsyJrA3UIMag2tSfd1EGMgwIT0whWeYm9X3zSfxNrQCMXliwcI+0fxDl2QgRICsBA5vt1tIffj
gSErR7EHWGEdIaxNn7sVHkuRc6oN1B4YNHBETRZcoCyTxsSzSmlcZpO5AqGgZZf/UltK6yxKSrEa
xEX5Cg1Vpww2CvnJLfkCB6MoTEZE//ndQ6lCflm9NPAQ/vUbJaOq9T+IyV90oYZeMNG17P+hafXt
vbgG00gt8f06tsCaR87ookQ243pMAavSTxXMjDMnp3gGfZuNNu0ZlsPWnWxHOB/EcS7eTOfd4z1g
Ed5rOQSiu9qWqekRUSDy7DFEAfUGOmbAuMudLTe90EHbBlXLdQlvkPl5RmMqnmeEyGIXBctufuL1
MwNAtMFAbuznzg8X+bDHyaXsqt38iKwKUsmHeFYjy0k873BQrkI32Ef/4eVGLfuK9dfkLRXhXdmV
amgxbpWXHC9nmPxmFcObXDCgh/hKuAhOnY0GcXID9HlanwnGIElfZja6p672QprQWLokfbgPXX4k
Df12BDX7tG57pgHzVJ3+GfHiu5B2j5hdblEzqGcIlv2G+asZ3KmfLSd+HYuC/ziIjziQy3Rxnfyr
ZPHA58zTqgGTip0VnbzOZV1m42m1aFCHEULTcp+PmLOX2jBiEDUTnROa3JHzu3kLVavtJZSFPdU/
J3aLSJXcYX3rBSb1GtYpjL4oCoawm4c/xD5yQPjeAM4YwaJpyAQJhscjBc6cmEFJCBRpI0zA+Tfy
C4GIVXT6MdauhSaaKCgkuwq5Vckf8fVRqukeRYwpEJXd4GRpqyioIo7TpzI0sYcHlwxyEy9TlmrA
rpgH94ZdANAKLI36D4Yw7ehOs5lF4efO8lmt/OwnnYx9QFhdeoCtYKQXUwgUwxua2cIgelz38MNi
i1+TT9IzOJQurYjCXyoXWOW9VDk+vTQf1V13UuZgOd7Z32QeUFuVSQHDn/gB+5VXnBQ6K7xULF+F
aOCIDxl4bmyiq0Ha1w+wK3XV9PAAoEiVwM8sICU6Z+u0LRQ5eyapKnmr/pBUqeWUFftE3nzsNSP9
Fu7RluZbSkDiXFH/uox8TtahAqWu/qlaAdbcYzSX3Y0ndzzloO2Xqj9cRyg/rCN+AQWCKEEh5Q+x
S+hG6bou0r//YqxE4Kr97s3WZJ9LygSp0yOqRL0v53EF/60w/os3PaRU0zILcs2ZaL37aUeAsy96
wPDWv7TJ0D5pNQMDzqjhcyhJ0ZVrAPkDf7qEC/aH6lm0KUivlsX9TEkxkrsHyxNzwz0DZ42pBB8e
WSatenLgLlEtgCB1oFoi871dpVRW0Wj1WQs8XihaO2Dyxx3THqlIj293Gi9qzPvATw/TzHbJqIBl
JkeztYJ2s2IEp6vgXSkiY64ckgRAAFdbajCebG0WJ1AOqYcJJGSXuCfpL4oZJUD89Nf/7uzQm+Q3
NlpjEudWRbE+0/hejSqV149hgIeGC8qR0LbE9qFHxh29wUhcnm85ttTkkMCgCNL1J5jmOdLC04xt
Nymgb2UNjTgIEjhooPAOn+UQMFBDiaH+69h+LYaLkGnlFdoUUYI+DURcFnL91YEjAw/W9tizM/vu
R5wSxs9OH5ocqCJJe4DI5aMSPz9ss1dTLBuggqXqHEg4jLtG/XnQlOhEGQQ6hZMB8v5LfmzI1S5J
xN/hBW/SOIVRoSdfFRzKvAuZgpVD2jRZpTLpp5i6aW3ozEfjmJ0YYnjIUvepAVZvzq2EciBjjRgj
oVE5h/ATSIn7pQkWHfnwcUxzTa1t2pyuxiY1p2l4BRHHw7Mve1tsSpnl2uV+EWawD5RHIkqSycAE
BZq5c7h0ldzPsBWxvOr4a49hAqU7iUYshc3jsZ8R1mZGH9GMNP+kdZNeArM/myQ+A3KnRJKznPN1
F8pbPRsY4+yLwLtHof3VOCM7QGVoq6JQgW8Y6RhmoJgJTujfY+SFu2eAdGGT97WY35cXNDssIGzd
jz5be3LJeYPIljVMZQvTbdfcqaP+3leMwRC0ChimuYqgrTiQPwfy8WVt6efscbC58u6KhSRCyKXz
rNece0S+XH+Rz1goNwxntYn4jK81o3p0u6qD77XqN/XJk/X/66/PzlnHI4WINYsiuAl2MH4rqlcm
zBOAvtTbR8ElL9VlR7El0VAJGrBo7RhpSgYGp8UueIzIn4N/fmzlyqLuesTVH/U5am26M04P8VQd
dYl2lEmCHzUeBxAZO+6tIyPsKiME3mtTuO1NEwRiuFlpaht5G9mBybRWVUhZSQYXaK6tMbvjjvV/
8+GkoolaLPzwN2CPzL9XVtU7woJ928irwK+dlqHvqFF+0ozYmjWCoUSeXFNrPDlcqrwx8Ghvtnhc
xqaBAF7u3fvzKulbwnOiA6x6Bkd8GeezA/SBTbt7RKilprPith9wIf7GZK/hGaonG5oIzP4hoJdh
NLR9SOn4anotlritksbdCMEDzhv0qna0M/XxfgsaNZ8mpWUsm4u+WXDjbxLB/8/q9g+iaRmrf1xk
1AmTkx+xS3CIjE2tsvd44aQhtK3MNDSLEljpoHZVD52wL8RWEU2tRVDcu6wSjG76QzU/kvNDe2lC
l0ct1F/W2VVIdYaC8WGKP2nWlb5nb4XSivKF0w1OwRv/h8j+/gVxTyDXKbb0kysfqXFRnps5H8U0
BuGK+eeEAjVg+hnCJJ0pRlcGPJsmVHjVBKff7ShjBo/tjcDoTDup/h/83KAzO87DOKkzzH6JMghy
0eG8a/BnSHQPNoJfLL9Lu3+dcGEFDJTwZGjVV4GMu8/ZfeGVfTyoSq2Rt01KwEXMJ5fOt+QL2cWB
RHG82U0iVb5RAhhfOHPYZcQm39W/ah5mBHV6E+0gcuVpMBZQJss2be/nPF+nMx0xzrOCAJjKQ6I2
pXHf6GrndZKLaE6H5zjtygRWA/b2duntoWEg+1Z41exz/rcKrXagNXge7N6ngBbE+mwh/OnfnfXy
TOZ++aRn+pL73Hxq0VRbLJgzTIzVyOAWa312GJ/XJ8qtSG0FbN563cZ+QFM1poXTe2m3Jkk3L2xD
bkp+IoWmE5iaaCT9l/HaHkfdtLGkz/rT++iXa23+G3qDQoRQ5J+G0UdyglP/HkQNg4zC33AnQUkZ
RvCR5raAUjmVFbIxKAxtg+jZahNQYt3+iORxz/fANl7WrpmS8EldXv3CssTY0Rw5eTPgKM+cdHjb
VQCse4XbFOYhQDZ6S5SucviO6xgJaKxt0fGpdseHnRUidaNHG1xsJ/WzPxVItexFzASEljBx2ARd
KUYAck9DYNLFjyPwak4Iad7wHPaUdT4UcGNWb6piNWguYpqygpD7HX9eE/Kh5pIWVoOuV6iHMOJ7
lXxMAyHOOplLfqdiek88AUqi5GsyNKiFabmkUl3zn0lAy9Ne9guNQBEOaluRhuuIZCbiVU8NZk1K
ErDAUpHRfRD40nHXpV9I+WXCBpTMps80R59gqKDQvaP0ZdKyQc5vVftFtVuWwedU3S2D5VkhZj5i
pHUpgNm1IoXbjvvh98lebAZPorZDYmZXp2ihSpYU/P5Wu4silePYvaaR0hPhwS2UO6BaAiyEdy0V
E90mHV4xJq2yzQ7kzPXDYBC4RFvhYhbym3RW05+HRYQ3PlDE4RzpYM/09hmDG877Um7ZI+eBBrmZ
OO0OjDrWV39VoxhXyuBCTqBS79p8XLTBkcvmtWVBMFJe6yvZLN7CCvu+O8OcoC2bAKjvAkLCScuL
arP/pZ9yVY+vdOK6W/luzu+IxPutf87ude6lMUKdErq7szNBJB8W7R0sAbHP30ihSKAYpqRGAM8B
Y9SaSGw+hUUhd7xX9UuHSpdy7YAw9eAMbykGr8ctBP7m/c2eRpvUDVtTzMMZHrgGgDvaCWpjEuOi
89XNW7Kur9UJHiGDe5z1LEJGcQmeclOSlNn9uRWOA1ZS1Gj563KGCyEF0XLO0veuYMPeuQdobbLW
NZrwdKeaHhrAKfJmCQFnxrAmK1dsUusOFhTrBPqSGxYcAdGp9uVEqyseYwvRTUcYpmApGw1zZ97B
EZzm3n77ziKhl8j2iU+FnPPFryOcFNLLlVrQE01rYpKCNcf14TAq41T4lZp/XbW6BQn1xZD7MTzj
ufxjR/sTu9YKBppw4TtWcBDZJawLOro4ktBTNamHQLKnEFRcjOfal5pJY6asE7S5kIsyqYed8LXB
qpvgJcY3nWfRzpKqF1HJd+qKn74+9pBdhKhtwbyyG+XHrhrv6GQwY13rwYfbUg9QforJ6VbIxU/z
Fb7YKNzNURzZXdX/quky+Bza4sIVOliWooxaKJjWZ/EAGRiFdlA1/ybjBbsjo7CXh0xxsWa3IVqm
cg3bFVUvkkx62czG8KMrrppwHIZDWKeIRAS85QOA70GNVU/Mbo6kYm6nXANBB/uFwtKh8xuY5eLZ
E0jhJ0Gzf/uXQ3vfmRs9bXcDhN/TCEyoR5owqWiGE3gxOwxOk0VEmkwe9HRvKfaQ+PLuVPoXh8ia
9b17VzYprUNfATLlqKRm6/h3/qylemjebshGymly7dJ2bP0y6XMmk2QNSekiCs85xAMIhStjtoZh
K3OZtmVVZ97tcYF8UlJ0oADxhlpZkugtjQQAUIUdw5g+lpSM9sx4IbnwqeoK+kI2a6tFHOsrWtRe
9sqm893aAwFHecoThoqSTD3n9a0H8ygWw02YTVJwDo7BT3laFBotJkK8KRhmsGkwtWUOkfI7hZEg
nfqBI2ycgrkR4k1bCSSZOwtpELsuVHeL05W6tl6MTJD522u4+BOfO1zjKsHhKogETUPO2Pbjsqt+
uYyKswRzDuO1BvaEREFiX4K7y9p2kaHLskUrzJMpH2u/LSfZHy3AEJXI8GRVayPYkjPycTZZ2u8x
zDM7y4/tIJv0yJ8nUFI2vPLb7lk8Uxf+uAb/Ml2baGHDWH9UKN3iHLTMEqw08rF+wEopk5VZ2WD4
vq14h9GF9aIGzEi7XRWnP5dU+cv/5keLCahYeE4jY+06kr4m4B5Tz64KPjLg2m1VSQNJ2+rsCD/9
zA/veXxR137BQylptjXWCZbpUN8C+dv85zkl92jrDbEW7R7/3OCtPYBF1LPlqIUH2b/TWQtSGoB1
YznyKnXzUcXIr3Sq1agvx7gUa8JPzUNFtY2ZHU0xGX3C/v2ZbdLLaQIZXWPEvYWt2TS7fhw/CnuQ
2PiSHpCje6b/ZRnYe1+zjtYz/nLCoyE9q5lNG1iNaI9sLNojWVrVamINV3uiubvwBjKtyM96mG2x
ncvDnR/I4FRccjjMluXH3ODWtYROyZWyTdrsPC+vGy7rNv3OvAhqjGEvQ1kKb+g+3aadXjMR3ASe
gyQoygBrHi2Q08E58l2PpqmgCnZQsfdn1lrqpHHcDaC6rMT2kdMGMOTYNmHy26e7PVcMaUeCHS4B
BxD3XXOG0MTbbqQsNztnbIOEdiV132FQrhHsDTgqMqBsN2RWaA4nE+6whkJ5hxbuPe1lSF9Pol8J
lD08z+ZDK9cxqIj+XoQnyLbGAZU/fBYuVddft2X9s6Ix63NBXSloARr5ClCLNYejuXuS4HXY76Q8
qfE2r5kLKzj5MLkzMot7hVgrURXyWgUzzcpvB9R8j3uR9RCDE/nnE1ZCbXICh6hC4I01JVFW2hd7
MmG6raWchJvb9/U8TDtOhq+R5TCUf8hSCB9mjFrz9t03p1YtiLB9xy9oxqrWyX1se+tzfeWHfMON
yPFK9Pv5M9sGSOoCtrSPMAkMrY6a6GT2SSr1ponx5DhcW9dZWwJFoaX+LcEWXX2diIle1VhGlc62
vM0vGG25sJJk3dewKfqUK+zGeyq8mnEL6PYkY0tpUAb3Gh4ma++Hd22oxcw7F8+IgIX6ZWZGV3EM
7gVK1yd/wsIf3Q0nqX2t1iSl7prwZpbQ9EdEsMZQMrbftYMl26AClxQ3F/U4U9eyHANgTsi3xu02
qE5IIfsYMUITlzGPy6Qg1VhoJNJvr0tYS9wutmoz4u/6XGcyJoBwttfFiKXwFxD12APVGhsxNYOo
9FDj9QX+aGMdF92sYaS2leIbqKv9i8CM0JPjmaW4+pR7a4c7MvCYBuyV3o0LliLAfxfAZ0Ya8vj2
oizugE2FgfmttQOYqwht3omwPFImWUckNzbRvN//3K24RqDlynpFEqCT0R+1XlyF4Kf+qDqQm+da
oBfFQRgjOSwc60S3gpDHjemWBZXvM196/PjC9aFI99a1jF1OKd/gOeYnudEqedMvdaI4YvhthN2h
EbC0TPA5DOSOnGwrmTFBH1SlhYoGp7KwnaRfEYhkZOJMjbH03zCAJnr9flcu1P7WkzGs8jjpg58C
0+3Cw6GmXe1CP+tXpe3rLRehjlzjYYHD3ox4EO7Su3Pe9cGNFUYacywr/Zty2n6NGF+Jje1blPeH
77OfwfDy13Uz/q9o6S98Zs7OMSdtiBjYWTTWI47TzD0Cl7pW8h1Nwl/9H/pobncLDtB4kY9N3/QR
ndCtSNbXygjxzyMvtfhaSLPV5h5P2G/wYhIGlWKo1vi+8sDC7qfZ12XfnPEqY6vI6Z5AB+qQwrGK
7uzypIW9DEyaW3TKExq3jVALDOsxfI3Y3U0zFCohYpy4QQVXEJP2pjUPed46fF+iNuOhEbD8iDHC
56bIDotziG+TLNlS8I1x8LmeB0y5IWn+HEKhEXnMn9FORx35r9EmPi63V/SkDtIJAMR6FIFKYxEH
YYyrlFSosmPMsIQuCXX71s58kG8gIANe5e9EGNZU4YX1AQHYBGNG1/kZeHzmj66Q5lXyMPxgAElb
5w1adydWZBY/JWPlttdV6+r5qmsm3wz8Zd8ejMApAym8UU30CoMNmYWNl8lqaUbIQPVxo8QnuI7i
svQf75XKEM2lF6uJSAk4HuEjDv9pW9udoUflgWpEAmfTTb6h0g7+V8zicLjRrLL2o4eSHyt0OVNX
RvuXHOj665CvJGU/3z37JJbooKuEZ7GPWhPO6yhvDmVLvOg6fUpLgVLfAmy0AYJVk39djwERg9Po
BOnex56dWNyhFPlcgq+LCoB1XnPa6vBDXu8xurJw9VTFZ1jy46fjXPSt33lP4hyFtgRuKz7qtFzI
oLyDvTB43A7BJUJhb/KYnUba95FdtWazOwH6dWjbTt7OO4ZO0f64sFH5U5lklOor+VJChQ/sdAMr
aJtQ1qIu7lrX7yDRAUXs7ORQQrBOVFBRrOfbHPv5i5joDKU1zYmRqBPZcuAkWD0wXqv7s+9/fzWA
Q7laTOBO8GOYdQt0dffGbkfuHxKCBdo56rF02dd/N1zP4Nl+ERNMJH38VGbsQrVMeAnJlXgSB8ly
H6BICcHnSQfMLW7Tpy/Qf9cutS+3gSyZCXG33ygQv6D56dFIzcYDgXOm9MRMWVCMe/GORjFptBhZ
zdqrPHXsg3cFGUWk5yMc8dfh4ofbYSWZ7XcNZDCAQQhh6zeEzigyGKcJKIoKjR5CnToXAm7azfwW
IwGli1E6W/YOarcoB8f1G6NOTRBxbTEP1tr6nXqJCP4E7o49SaeUhyCSVept/qDismggL0+HQsAs
vKEFAQuCquyHiCq0rE9q1St0t0EFrP7aFh44e5fZFiEF0IlrDtUG72ypuIweGADOmN3GecZMM918
2Q/tt9gFWXflabe4uVf6X8C6QJgrbsN1m8bxNGypb7M9avjvfUTLpR2SDE9K8+e+CzpZshfXXtUi
gbyHi4bmwEWbZWbiv76Fn6Dmaatae5P+XPic+zN4HJ6Ha9hiqqNziyRpApNVYAqywh3hTJZCwHpb
l+q1n+F+PvJvsHXkJCO1NtfwrrtH7r/Q532tfzDLmlRaMN2R0SyDA/OMvSfo7/WVXbnBobP9ODTC
BeNDk6/Yg3bzdTuVBdMd5HUqxjCUNpo8d1+nd1AbVgIMgBqyP5AoPNpfbxDw7U/5QIfq+ORLS+Ve
cr5pgjOkMsf0/0d0sHKyFRUKjpQwZ3dyyIy4mwE3AwaknJ6jBBnveqlGxwbo+FpYdEhLrk3NIsxZ
Yl/HrcLjmou3zrgWZwehqOwakxBYWAnSxERCbfthIq/PhsuXFX9S4pSQvs7KzZaUXPqtJFZ9vGVr
jKD1BjGe0iTilkMkark135NjhAPsQJg/gAVWCjLxSWCzgSJUjsvQsDj/1xD0WmzeHToBal5jrWUb
DxOmy0tEEBPpcN86fvND6ly+30zmHvjAmPn1WzpcTBZ0KK9cJDtr9vZpjV/bWpwWAsqtrfVUCVEx
FxHywlQmryQbMWBXgtcffcr9kck4A4kSFUSgMuLWLCx5Fg5tPojQ0Tve+ySZunawjdvf8gRIHnOI
YIJt2FhPVd6VlikrLsTrFm/B7O1+laJYGugCWP2BJxvmVaOSYcG0Gf5twncYipUxrvsX7wELTTDg
7u09DX4fk3n9sza3jb1g1F/LNk81tHulj/vc5GgBTB4/wyZjJ8lmuJdgxeRiw492Uz7ym7Sw8G5R
TBJumL69z/VddmyAq+o+j0v8NoIbCkl7uTS7dnkJcP/a6cPwRLgeIfwEJJEnx6s7DzwskIQh9je7
hjfhohD1Mh5ANFNAmnW9ZrGFnRqqrlemXE9mTXPd6DrriA1FSH1oGQ4BW2NeG3QF+FvOoS8ihPcK
9E7H6t7FBH1GRM0Lod5R/g/ifAP2AnVwkNw5cbJ9g5N8Xgd0hn9GWbORQ1z+XdqGJTDJgW8fj0pR
m2jGFk3yIEPh1HSz5xc/KLWZmAn2G2NG4vkXmXrm7FmIJ54Lh0wyV1KK5Bl4ow8oq6OuxS1TsbyT
FIxLFuz3LSbuWlf5nLr41JrW8HDZTs+DtjF4VyAN/FuJMBym7VNpbeO0m8GDflYZkB0PRK/m9gCV
7ZyT2iERLXStkg8EZwkD26SLreiDcIM6/gDB4S5mYVSEzc0tmiWqcaKbQv2Bi8JhUHN8ia6o/RCB
0dyGsdiyo3Tc75jp3nIvOB8fOwGbbl6qnWY+84qe+9kAa1h8nYV/mpnQd/7jvQanNVHZQx5VOslg
IkqgMgEHJexODVy8UpV0DmBbeWVJ4ABxK1Mc+xiAU9EMhLMmIOtPL4P5bj1wf+H5eeQIrCHGROaY
d6pjGOAIEq20qdAcElKwkSXeS5gvEvGgEhvLB9mOKxtY6VHhx307ODCjQKMlubpfiAuPQvaDfd8p
fyiXzpiZv/ll20GgFAhT68tep0tJMBXWER07n88iQCzAtA7nFzUrexmhEtXG6LSvGDo25Wda2XiI
aIExpBJsBX3WX7aSmRjZpwwJBckALZ637xAATWOIO5p4+6ITDothDe5WxzwAmybS/IEv5xjpogBB
bInVys06OUUia7dSSo1HKPUJp8sUaN8ckzSelUz3tyUtxMYJ6HcMyVdhtI7e7+t5EseiQjsLRAsx
ZWnGb9HVGvUO4NibjDPRnXzVcwv3Zq5UmsRIOPjWdSmqYoj4VA+VcuGVcmFhbTCwpx0CyzIp8TXs
+atpMK8jTXT2tHHVdYP4F9oittqNrs189tpD+hKRjegY/88QZKFdIL6l90qxRlyEK7n50KpY3bVz
rX+vZDnh22Ka1v3MXa1UGXivDWinYC4ATIz5bwPLV73OGVBXfh0rWFAfQzti0sEjMRDwPZgzUkiv
0hyt7yZRW9QRwP7Ig0etQR1Hr8+IYWL1Amewp76nTRheTxCvXI1UT/ZOzjUQkRtuo1b/HNRnnqXL
bX1aUprS8TnQDsG75ldKEmLxZs0iNAt6PTUQi4TlH/iqWiFtzefkSyIRm4f9rqkCgr40ufeI6Ufo
w6O1ITtisegxhNB2N6ENdZ9AyFP2zGkrO4oQvKhElWBHYwdRlNqhsErat5sG+cBH3Q80CgUuDY4S
hSqMy+U9eYcSr6ZLVnaSqPMoagEZO2GwUkYUeh0CHwP6rRHouVrG1SMGjY9g0f5MjUwc1wmVwnY5
RyXpDJXXYDElnGEf5CUT3ayL0roNtxPpjfPSQrcNYDECDK5SbBnbByP8fzq3YNz+zXZJk+tWLvFs
XRApq0Ps14wMLzZUevIOsIZ51mfEdh4KpuLtsVBexjP4sIlstXNd0z6yXpRMwV10vG7y8pteMuPS
Ld0AkdDl2GhCF4oEg7a5o7DPLTyoHxf8Re1WF2ozqLe6vAHj1hFX3fN1lkpM464ndikByOePXoL7
qo5GNro03UZCUvD6IBx350gOAodHWoAHWcWF6GB982J1rtUoFvs29M0E4Ul/Eyxs5NezzhAJXHGs
Xyp5ua9J17AVLKD/6t3VDykxoVrGTVRyofidnuIRBkBf7NH43n9kp4xOSPhyOCJuxz0bJ5aKMbmb
sBWkRFAqekaR9uQLLnbr7Gj80lndSewqHTI0cRPyKdjqzcFp4eF4yyZMcAFZ2UPkAYHauIAUGj3K
GLBn1HrQi5QeeTbAs2i8mk5VHvY6nxyuqqar0E68mkCqWLrb6xlKJm6vCaZfc2U9pdhfMkV7mqwD
AMB2sp2IgGRwgcKqqtCN/crMszDHsgkgDk0kttH3y4LBAAhjmuHGkUxV4IKKKkYx9rJRnJVTq2rt
j8q5v9C84Siurl8tqX4xtaIvckRc1SPKTGNYVR03ozhqSS/FtLO02OAjkQKdbJ59vffUrddFKA/K
KbTJNwji/gzaH8XFp8TnoZudzcRMTYRza7sCNvGDUvzvkcnBSuM8nn+cr+W/h0yPb04uyvNVnaep
BGVeEb8jCIFMYx+f+WyOqKk66LPaImCpyVvZE8U92Oe/AIKtL2xYlKgBhfY62uwup9wty2h86HtD
vLOl0pKhWBLD97e8ivBeJg0kBv9oOuXbc9znmP2YafTN2+SvSvtY0IvIrMHY9bQ0i4Q2b6d+K9Kc
mHeYkO76F1LIlm1P3ypIZQZapR8St9cAap783MQdKMV2fYmD2JDRDVBebQ2KzZzRKJ092q0g14kF
KU9b7jlRM290z8qz5q1T35OG2y0SQDqdBzipgmSBJO3XvjEtUY8pagC04Y4IFj1jlxOz8oFgY0BF
CovOAGN2w8qfUU8qMx09VlXp5+dbTBBJHhRETkUsDqB1fMKHFEcKFV6CssSteGkcKEdGWDPMZ1Nj
TuqarXNIZQJ701Rsp+bsBLVCzLFkr+3oPBVjpQzzom3HpOUa4XxVskIZvs9l8Zxo7tTs3cpxRB++
YXqm3R+5Wc6w2JmeRltskX0sOV2q4WyEhzwEJuljK+ZmJ4uCBQd0ls2fy2ug3WpWRGRpYtLPO7LG
U1xjUtIc3svkeK6Cn59+N9Qh5ol9Kzr0cNreMQ17Fg/Ac41NX0/D9pbwMTzqJF5zhw6reSWAHBHy
AjYpry5x3Wi7VzKMGhqCUswOV//ciY7WuqpAF7CNsQoheKH0LjnqTijLANVpIW6zygix6gbXMtZu
mTx8AnRwlNbVeSWlnZIiMK2UVdyNHUaLL94yFs+rtuOI8i41VlX9w+UEnoArVHTCFvrzikKQXSk+
LfGO1xe5kRqMFP1xTwdfmIoXdHv+oIwEzUd0aQL2Y4obYGjAtKIThPn5CTrMJJxxcqo2ldxWeENK
idSQEGKxcLVDmq4+kG08m5QgNcxQeoi+w8Em0G56/228UEMJTbkzvwgZA41Gfy3t69swFMJmwx7x
PnONMvlhxE4d/ypWUI7gRH5mU3FFRmEJRUedPSXQjBvqiyLzqii5SX1GdGk2/6jZ37EFuwF8iaos
LIds/NrlRMLpI4JduRW2GcRmMGi7alWyWVPPWJDIaKzLmoFFlv5T0hBBUImM7gYe0Hv4p5TvU87a
bfSjF/iycbiF/mQXRqzb1QasekulxUCbWYRl1rIBBIs0j5eFPJk+gCCbcE5fJi8oZV/xgKQ4LIgO
apxod3AuYnzCiFEt1wmM1Y9JXKg2Nf3rASSq5yp2GunItJa+9fC3EiCvo/8lNj/mT2jVdIZqhDh1
yS2EaLHD5EPD/HL6gvhQKS/SmnnrpiaQaiAhUHF3PlRGXvG7JUIY3bRebAaI2ra5vwzdFkHl98tl
Up0PSp8ZpTYs1yHq9+fF6sHOutIJ1037mkfeB3AXi5QX7cFUk7cOLbmB/ks2cnZ5RiyWAk567M5k
tO+dCnXBVNxUV/TfhfQg0mVTkqqzv6fTpDx5BR7kKy7jYskywXumhaTM+K4xAgsLei8PRKsgx+ox
XIMg4AL2SW04dp0/uLPm0M+NCa03NMZ4izdGQn0qv0LcOh1H+8+7ICIygEiYrk6f3EwQApnOQLiG
KxY96ZDqrHFCz+V3v6dQAD59UzcSBwDskz7gAoQAEk/oXDb/KrA8aZWd7EjnK3H2Bqhd7pZzYMTd
BUnGt6prk81hfFQJTmMlT1I1AUVQQd3Wdohnmyyb8TgWVrRReLLotf/XRQ0YMd6TPMcDeUDWxb/U
kMfy+a7Uxa+6QIm24eonwi+zQLKoEGAB/jab2VxQf29Md3Mf70V3vYoUuIEL9DA/OSDDfA72v5ih
xZKPb12VdYBqJQxhhZPjhD4M7VhEmNeVYGjrbMviwe95trxrd5SpGSeljtFEOBG1j0NQbmNzvmNR
EKD6L4UgKHa2LNOIO8eDjsG+tKo6ScofQg+xmK8Mtd5fx9GGpV6Zi7bSAUIMPvE7Sz7h82L1pv5S
/Xk+z1jF/gtXF+FFLF6inthduVZQBUc1Q0nXzfgYYV4qd3hIdG0jtKVy8UZxS7U9V5dV3/COkDzh
N9j/+4OaP38Se+For3YMb74wdkWHk8Fl4lVfDToGL6KcZ0n1Z8h74g1N7Pt2AsosYLMZOYCZ5TAs
GUCnkhhC2IQBkBhQZtY/B9UF2HMIEfmoR88PlN7DgKg2xB4ip5AKXJbFipgH+jbe0XB10P/QjqJO
n45WjfQwzHU8uEFJr6B6RHDs3hXaYGh2LVxJLGaqdLBgrISAeOwfBU8Ois8OsGai6U7qWTpAs3Bb
JwAhRvEsFQlW8gKO9qEQbrmsAqvgyszgG3Zqj3SgjPpYKA7Csw1EzY3Bzs36AQHUFXX6QfAoZMJh
CuPC9lR196rkNJiGngA4MOIFECCBdRu9uC1vdG9YFtpLA7ggyA4x+cvrJ6SUBJ1AXct5BhbWBtnE
cOOgSc2jQcDWqbtky3txHwLBcuepoV2dVl8nSe0g4GXc/TzaIFLANUwf9IQNx11cDkeVSKlZtEBv
gj83a8D7QUiS5/tqgROBW3gPqSjl9yP/053Vt7Hb7R7dhp0SAAxkSq5Ebx+PTNbtKvf70xpsIzMS
PhkLHIBVN7WSCdFaO9XN1nabaGZddfhU1DOQyB3ikeV/a16VTGKwf2yvOM/8FaRKOS/MHLteT4kw
ngPw9ncyIkFjwWkAJb2ZgG0fxZQ+QUzEWtpIlUYoP75hEGr6NmxxOuIzKy6mTFFAaktWkPR7JpbA
sLtrCS/47gq07POHPsIPGcs4vMj5nv3malN0kGUAG9ww/iB96VPFmfiUtrJGDp4y9SSeXw8eAf/C
ztHb2jTvE/iPXRFggUEZtKUCkMuiU8jaPwpQ6EdoCHj/TkMkxkXN3unuy/cg/n+MBjD+hhFVSn52
2CbsiAF0xaRNmWgS1KZkmOVjta0AjftH8mndJDABQl9cYNb3+orWGUaHyslmaHWoAxQPhpFv5vqh
Ac5bpIA1eAQkJ6sl3+kjaO/fB0/uS493aIYQMXb26/FHz1pdrJnp3nXZhW2FbwVGpo1mjYHWaunK
NYrl/TNwEh946YHerYrJ5BozQcnOLFz3YWI1v00djSy4nz+Q7l0/16DxfHtjWJMieaWH/VrrZBBv
a7ip0IcyQkr0Sqln+YR9BhohmXd8V6zdEyHd5+UiYFyfhb/Tl8P9JrC2cbxDKiiZ7JXS1WiJUapw
DzDkPch3XnIltXwpoVlwB9kkDuYQjLWoyiPwgTYCXf2a8uoXmcKSSwk16sf1z1EN/iS4yan6FsGu
CLB/Lxgjbiqg4A0jrzw4IrVn6JTNfGlTXPmI7lKai/AYREkJAsm/ITRVFo+Mg3GEbG0DFXE2Abl4
rVlHBTXAKaOuB5Ref6FDl37cVopLEoiQ28wPfnsCSPxaf+ECUmmHa7AWdFxnjwnB6gaVVwgBuNC5
hOofSj/EoQbdnR8GStatOrnzBTliqozJ5hp3ORjgVGzJLEa04r7k9uCw0uiIghi1aqmr0ZG3kXLd
OzQwDK7Tbs+FjckGSccVmYP8lAs0LIcXOh0mANmOaHEvjq/U76/ecjZSEcAzNyGQC9OFGc5+swTU
J51+hFOgENfgrO0ann3DG41i8N+fXRuVddjN0FZ63Pr3pBK38lLMtbJIbDTdX5HYHcsVt+18XRNw
CMC93FyOgdIKGZdMcLwgSPJcg1iFU5+tGIhV5k2qe0f3fvZnISNJ9XuYKZ+etdbbf7VeDoBqTrX7
0q54OnBUvp2gpofEbNKMTJMSW52Bgk0P10FWtG7LP8vZAdJvpoAefEi8DRLAUMP8GKpDRIG8h+RQ
bSL0gafmYGIesKtkcioKUXNL9Y3EHqvh/7/BhMuaVQVO6KgwrrojbHPp1sfdklraS6WvlrE+M3d/
EMTqUCpLgTtKETOXwPzBk5UoRZsEbFJH0MvR5Vav7rxwdCLq+/AJp7qhLbew8I/Lff+jD3yL1wO7
csHzHfMeiLUwuReH4G6igs+ZqNfULtj3hRS5ICJlmgXqulYoreUU3P+BEdjk4lx3BVeuBetqr3lX
ds0EurLkgQth+HbYxwxkudN+5xVE92S6y5XioWebm1A38qVtaWNP6H29gquHTgXuxlgB+LuOFP2V
KkK4ky1TYrI0CnJxDS4d+ruZQEkFaC88HlyqQks/4AHGDFdPWY2XYyktgMVD6uyPaEiX++nmfong
PdUzGSr5+22NBDNh0dfRIDnlery0OZ1UaIg+RRD83yyNm2s8MQSKQ9fU6n6c0qkE+6/ZK7hEPWjY
TX9We68AogF3LKAv8ikYwxb2TMQ0CFh1foDUTbs/hzbczzY9uqwzkT78k4UpdlOrDCW5xeCUnhYW
EQMdqFJZ4jcN1xLUY5XIEdbCofDPtgZJJXRWXwYejWQH9wXjU4WJJI9Q62SLv5m8P/S+0zYTSVhZ
pP8mAI4kiy4C6H29PY1QvR69Re805JB9HffKP2nyzKUK/ZGa+jMBCJZkSeqnSLzRuk7ZfJPn+lI1
xRcAwX5xyz/Y3MFG1MxNFAbDsXAhAz9UnN3bIgRIjSxJI6KvLyEJ2SdXfLiU42HFaGKjZN85tk5d
6Vjei6W9Iyvqpmhucrv+L6AZXpniFMJMwrSRFWTEdBhvM03monK1wcpCSxL6y3R9LDjSZ+z0scx5
MHy2FK4EsNPZb6VSDCMrP1iTgakVMLLXBSeSMb8SXSRbfMfqKF1+Zk12rJREq/3vmz3WgH0fXRhf
ogo3Z50+OL2qWWFjODhF2x4pDS84T+GmTAJYVF3bFOs2QuahSdQ7Zx++LjlYWlTQAmLEntO0C5tB
7y0zieeIIbxCyPZt9yNL45l4S4T5Ef020CC9BDWZ4wdtVtIMFtXhqHElVd1wovDKvdqrLggY3mGH
ng18LTX0Ikm8EAgUP7UdLwIg0K0MbeV8rnpVBcm73nRYtf7yhyZaoERnvIXyTVGm2VVDgf1yiurm
fT3thpa6wXqwycfmpDdg8IUG1nF/2EfyodJosAnmPOxiDGBH0hjZMn/qyUUs9ODX2ridhNtKyrX/
fUpeII7uSHptpWNnx+PnR691QFPsqhUw2x359ze44OfbnYxtpDohYNGIHRO8dnm3Y4K4IWPg3V42
uyR4fQypXY5gPrUX+bxGD2zdee6sn9tw6u8auJ2DwusDIG1F5VtjUabnHgRFenCbehH+xgDiwyhJ
Px4R8UAIHvuKfDnL1Q54G9fjlVfkJRr9CszOdMKstFvfRNwX1iPxsePSWr4ZwLRN7Vx33q1SNCUH
7sVIOEJzNjWKPlGYFkj6LgEVCKEndxQ6IHbAxqv63nl5j8NQfi5q+YPlz0x3M9/HhQ9wJvXdEizc
RVOQMrimzaFY+zOv7b0544pBXrKAMxmHM8Mzle+NTDgti8WmtXthHnIvPidqwZLFE0/NoC6jfcOq
IuYOu2D7nwkS/QlsY2qu6O8qpyQJ5JQBO7RQAjYFm/IwXoW6QTC1A1SgzeuYGzaByjF+a6hgGV+H
es4XyqluoNeI+CUE9X3la9v9+RaRcsnz6ZIAdY8NbvFLWJdzuhYa4ABPxKywNNNVOsN+NDmvkodi
H7122F38GUt2jJmjZ6TwVNR1zw5y7VHdyOXBwUThS2Ohs3ARYrqv0j5tCWRymU4FOWzfc6gOyBQ4
TTN4jDnsnMimYdlbjvp9EGS8+PiLVx5IpplTpI9o/pNELxL0s1Phx9nOad2BNbF4iJFWr5iFtFf2
LKCoBiwew6xKH1A9PnStwA0UZdyj3daGe3tk//c9kWmR07OiO2v/qzTJ/JJUyoj7gNYIjK7tIqWq
57dcQ2TeMzL2M7F1SqXVF29OMitZV6pcBOnDxHLHB98dk/st1kVb9394dZ2hKvQFAksLGIyJwYsk
R2nebgIMpt3+dVIxRIF8Q2AjnBDK8u+9mO6m1Evnvc8ln0aYDHtbK3yVQj4ylIL59i9857oOUU5E
Gl9HNTOiYMcnwKK/bRgNgeDnjjv3RLQmhL1RkFUGZAIaDUpMwBgiVP/W2oEjPk7Af9TCVGWjcp/U
OYJrGtgTb34P9iDf6s4kqIKp/6NORM1qRrsTE/GcZJKQ7NqQevijAXoKxAMlRCGQdyG9nwSm07qA
5kakUzONj7rtPRySeWvU3xfije6r41KaxKbZO5XpMrrkpuMIp3woBVA7JVlEsJvEgcQYHbz4e5u2
QcfnJQg6WMzcvjFCP5wf/+WGsx5LrKP4DKGdHNCF9xswhp0vaa1t6A2qJd6gZ+TzIIC1L3eQO2ib
pUkkRXrIZ17TlNmHbrJXujzrhAlZUoIe4E4Y1KR31kQVYqGsVgkOhu8QTYD2g+5NJNUOrt6q7Qmm
fDbYoD8Ag8mXBIXExKjee6xb5AQ5UdqiAfLjq+0/pVOBe/yv7KBK4woqhz1vNtqycJ+fD3U2QRYr
RSIWDUk6FKY9Wz27QXor2M/wzTw+pWGMEDqqjO2Gfr1kPrBK++ZUIbHQ95Flh/+QPxIRbyRQfokp
vMn5b57yId3NgFGYUkoCF2LedvRZ+cf8/yz2hpWw858NlHSmExy9fqLIL78coCOb4141/rdqSui0
cXpqZ9Hkp7LIuYGVisl2UKdAedUnaCGmk3KoU9VtNbndtKzAsC8NulRTszXqTLt/tn4+ZXqVS2CZ
B+vIbye0FcHvPdMbD2mlJWP9S9cCRYbxix70giD1n9nTNFxxTvDBo8eRS8kWd6Frzl9Ml8qzOXSR
MgurE+7D9Ztt1gUd+dEJXpR6pVwmXC7T8h9ht0tk+eNJxxAGFi5wxoLPFPC0tWxH6GwE7+YrBGJ9
n9GtVegBxYfVlrNXll+hLD304JzjyBTkC7xVGEwtc3Opyo4gBnVS7rejeAEylqeHDtu3R7S2iUwH
3H0SqkXnSZ6eeZQgo1j/gKIDcGYTeqVPwrjS5KU3zQx67lMhgTcx9wt64d/igUyKnh7YB6z0g2FE
6M2LpS01zz1bbM81Eo0MSS6AQnwTta2NZDY0zjGLKzWlX/K0iT3RLh9fQvnJwMBioMcbtEX5VOwG
wK9dp6VxvTh52EoQRckDEv6E4qWZWP89nqBMoTK9YxrTz6thcs2nlnesQSIc3eQVk0vfHJ0DCVUr
SbBwTU9+hKgkQ7u7zqYxbjVIxCnkZ53lzd8eORAL19f/P5jJMskb5z/rvMFXZRB25B8tb7P8eKEd
UirwcCxY0qiYNL9YsfYF+Sfv1doYV2EmH7Pcm7hpHnJeE8cNTf28rjhZiStJHKcJLAhPteIBPmKW
q5UagDFWaZng/OxsRt+1wDcFASUHEJgyDWxsJ3PZEBrbxKAUAE4lIqBpe49cdD6G+RaCbPUMJUgE
GN6ngiTS0wPcEMo790njz7C09yWIRFDlgY5FLuNmbn9B9DF+fmRQjY7Kz6TwwHWl1ZohKlscMDTj
Gi4Avw/rs2TNfEgj5+5cZPKprSNacY8cbRRd9QLdKSgMQMJFzpdSAsxvRqz+wlzVwrHmPl2ZWOXo
8r+nbkk8sJeviaw0bopLrVQ3blWJOVkIAUfewr/EEN/PbtzpWkCGGGAEByA91vvoDzfd5eA8ENm/
I1LOsnSkr1m2+czsusxQfudu6UaiNPMArviCxxB8phMvV6vvk99k8KbR12xGyHmezBX1O70UYood
hNSXSOFSO8YRBxl4mhP1RZC3rCm9jH0evaV5/Tb+OhisrzJ97gJIePNizV3DpSO4p2XePZBkBA+d
b6IFuMci7HggWkYgACK8ORTI4fQZ+6GFvZ+Di+78Psn7xr3hxbnYXHhHG6mG0ZYcNy4Pwd0sjckg
YDZRIGkNkTpchc6OQLzJM+7tTbJ/rrDE4py0lJZeyiGzhO5c+9gKfEktC+Lx81h8HH+u1XxKjk+J
Qep+XkG+VGJ5OYnc9LeYXVRLu2fzoSAI2QMGkXYWhOlFa3bITqZ9SxW9r/ICV73E5zGz+OQ1ZgzD
02rfEYLlwtnb4CLesnFXTdUSAah3xNL1pauouUUxDLkOjc3r6QaqHQl/mMNmHuOX3ZHqXUwcBsT8
Si7JMFCMFZaI8ab0z3gUcU9JPy9V4KKd5Jl8EaB3Wfu/k7C8jZM+MsbwyoqbfLTgNwkTxcAPyYF/
LpayAolYwZmZJZLfb+T1Tp+41PJ0N8EemqufrwS3esf8IitvCRT+XTTgaT6+CoG+H2DH5LiYDsXk
ll1Nu8NRqFwkoirZ/P7af2KZor8pva7iEJN+L4DEK6ivWRIuqYGAvvAlmrzWO8ezKu1PNAzcoo5I
EycxjYHxup5p7symqcjN80vut5RZioUo2dz0PXXy9hwAob6DRfOvPSujnL9P9+95xOJL2h+XpzDx
XUiz1j4YLu9H8nLTKUY6bKftlkslc4OZj1OEbnXNBUQilzJ6H9mJzLoCsRtMppZAD//uxTdpH4bF
kKI34YJI852RuzgzUf4+/vndVumfrBpCmD9UsXC/w+JzZPyWH/m638SRqm46oeq5+a4CH2wwlOp1
CpU0gVI/KY72rwCQ98hmT9QGW5YT8H5CBMgG2EUhSn28Iwn8WS3Qg8mLahronSq0CxMQZsCvn5Cn
CfN9yVBdpMxX01sqnteXISmOfJWhJO5AM8vtZAhshPHCcJX1SvX57cJD9/YegmXiRv99hGxvHs7o
fGhLTbBe/Sqjwl9MeJ8qARlMlLC9S7cGv6es1hFiHtvXh26ELqBv5ztqCKYefurgMyMm3iWQTxgy
WA67vJZBmg6w4520QLiXbdgndm3hiWmh0hx+Zuv0sGs0X3h2+CpQq7h4dk3+OKvjQ7W6PAelvfHl
TTH/dTPjcXDhEvWIu3fX8bqC8XmnoJf8eyULEOafqDgdExcjyKvAbwJ9d9C1lyzwSZPwpJTy5w7H
LSUGo4JL6HUs8L6aSM7owep2yR4LqPrkd7whj18dsBpGe3dVMvPUbc+Ady7qqz56K2bd8ezSVVse
PX5AHeY7QtryRuQ4QtfIirLnA9drsHBC1nOKNfletZPWrDapxaAOyFLlchvDYx+gAYjDyZciIdlX
VhtWfJS9iVtYGYy6VwLf7ZH1R/sGNElUorNwC/cmHc8PpiTi9YbMpHtT639qUIul+7rG2mM2aPPF
BaWHRrGXC03wC/KxwkUgCVKbYlnQH2z33rAqiZotc1d9UteqzuYjbMpEV/UbPWiS5hqxy8uJ8zOR
Yke8Y3BC3XzufLsESkSQnSSqAD9UfliT9U4MbK36qKGSToyY5sXckHXJVCfHMjD8N+XxMntFm2Mj
lTtzM1E985U3A/gSBBrr9viD+ab67pWbjtOcP6nylvzL5vxyLYbgzoZrdnQeW4QkEy4PAMyd6ENO
U2FeSvw0te4KM+vDyqHg00d2DVWVQK6F2Fl2PSmelHRuXDueXi8+Mdq7psvv7MDZovJ2AFy6y9m9
aPM2XEUWs9/BNCcJweJhQA5bdOdwr5qUKDM8cTrtN5XAdV0NM6HIl7X7I7/j09GEem3vEaJxT13E
hnqce3jT0fWubFgrTP3cfKw4XIBQA3O9zp2xxWI74gjXdE8jmZIRLRT9duibsi0pJDLw2iwtCk9i
Uvh6RSTGZaaCEyd7A9fh5Ezcq//d7Yw9sGo7qPVriSfk2l479fchds7E7GnCiACxQTFqY00P1mto
1XuzXfpVSr5OVjJmeY+t4kwAsvL/n2Dt84GbO0DWhK6qixzoPRVECCzNWbe4ssCRRt35mS3R2MWJ
18Z99cc85f0GEwbnXpeRoeL1fJjc6BjgZk2RwwBKTeBbkFS7C7PHbkEEPsUDsnwhP7SCrfpSYbNb
fwHXXvmiZAButZwEfY7pDaRWxBCcHVQlkzhRNmG9dsaWSbVK03msrfvkU7QpTIdWy5qkQXb9oGhd
J9JaBTX7Qvn21KIaZjAhDmESswRLTk5ozJOidP7C0Q/SdPH0+PrPGWrZ9QFwv/32doNMbLqGsVgS
VGGIaVsuFZkPVfRztBE/ZZpfwf8QBrPvxzgZwgF1/gMBgTttWgp3vxFjws3lY6RR3nZwkUs4z+0M
MOQ6Tpx55/Hlifg131UGAM2A2y1/GxAqjtYtuAjQA7FYb5Es2oQpyvUI3XrcGQv692ElLIC2M9WR
47r8M6NJBmdbH10yhU/pDrEEVt4O+PVJEhzTVWudxyQarWiaJEGypP8+yv5vgpNTeIUYmTCzZhvz
yP5rwifPyaUd3l/nyCS73vbesxezAKf/56HevzeTO4Wy8E0+HLMXrCRrurg6drArgXJGppUecjYq
q1p2ZvD+sN9GDYy4szarHI++Wz/qcggKHaYFWEC+iZwy0IIJ8zHvqhTFaNDpAN7lDLOgoDSjGxE2
gFL5g+V1wAgvNICcrfVV50B//ZC38jU33LbHOyihu5uDoVWw7QbH2qFIv5j83qYgDDL5qPOup0PJ
ZtQLLNovj3bHnU4PmVQ2RkNKDi+7iuAwF04xDREaUIe98kdrYLWndihF+UdowKePL/ABUG+E89pL
W0U4T+fb2d5G3aPNE2jJhjOw8m183ArZW/jN2G6lMfs2Ww6vivm3a2kPOeHLBBivxKg9AKWIRkvo
D3ARdfVt2YoW+ed/7oOckfqxH3tOR4xZbisTuklzUsjLF5fr+j2+q4w/vbnTW/CSCo0MxUxwZmXk
f4r/Mo8fWTYeQH/9yGihfZF02cGvzUimOWeO3XzCnkVqna75MOgZtDWzovnBEEGb4viEdtZKwdo/
+4Ys96Y47T3oGWkFk1WEj2nvJ8VXEcd8RAoEcdYGSlsffI6aVIeO16m2o02828UsMzFgeD8n6E73
4lZxmdkgFcvtyLg8sL7yB5Yq0xV4xbkv8XuNxJOvL4t77uJ9wYafydffouwDO0Sf+oa+kbQo/GxF
o+K0Sa8elTDjwCX+nbb8LAd+OYhKCrCUznKMs3PS+RC9dT7udYwfZiA5FGYYljiTcFFdHjiwp67l
j0MSG3HPyKcd7cpm5csWzP3T69bKJAU2hKyeFJM1wDmhHNqY0hQMYer6IRenKGiz7DR1b1VyY9g5
Ez2yInwcBNYb4ZGSuwZCMDDnRKIf5T6FL1PfDEFyZejApjoaWJ7WLKX4v9Q23ZkTwRR7AmnomUVm
CoLr8ikzH38azJH6bDgvVjCaNl6BQ+f5PJCRNeT8RoWygJOr4VDb2SNpgv68aHNzVAMZYIeX3BaV
nw7aSTcUg0OhHJbzLruNLr7bN1dm633qC1n6HJELQ62Yd+oIZsgtUa7IH83u5gAqtG9r0bUOM2X8
f9A2Qic8dN+g02qwOnv91dwU9tIaKWysVIBOVFYGPJx8sHlFnSF+WQ4ENK5PbNu3ubyVtt6bu9z9
LBTeQd4k0NyAsvVUmsB4fABTLNnNUPOxJV2l0Ed7DqBQsCZQvWD51VwDEOoPJxasGzGLr9+tIr+C
X4oHNTiFylmXLcPSqU99pOk5K62YRZpfbl3hUZVCVvmcV3Q5GnpVt+a3qLbSByvTfXK7bBzQmuEB
bRVozh+TiVM485w0Zcb8plVoi/H7ol0dx4qAhEEYZ/29LgalYdT4ki5PMEMqLQkOsMfbzQ8AaTyz
1vfPs/wOaZvaeoI2Op1Ps+Ac7QZLUHYtq2sOi1V0HOqi0sri2yihgXqK0TKgdVcb+JH/HiwAHIQL
Sh2H/UQFJAaY3p9XdXSAUsvy37rc6TSUj6LZeU8SkA4W1b3/JBXONauB1ryTY6R1ZyAhdimK4NFQ
K+Y4SH5khyUhxq++MBowntlSD74pOHVSBRqz2t4Dg8bOBebHe4+13CvfSC+0bLRo7QxFSODZIi2t
CkMORcv2FV1EJJQe0uB94NVtxie3CIOhsnQE5a4UUvEvBTx13i4N0Toc0ToV5+bg9CCnoXqX4tDj
/aG+czQB/hgwBj0SFnYl/QVYquqiuIcK2lcTKKTVuES5rSOWQahbNcUxDzAGF7HWC9NFL+20sAM3
gHL1kjuBoJzVEFwb/Q8Ghjdy1tIpH6cUqCB4rpCGSFGzq+yKYhlpdh8imtU8myeL5myzRkQrugwW
JCcvCfDtaD+BkUxI05BW3av9riQ6EMZ9p1e6Lc9gLhwBHO9hF2utK/PeJ5y4LgYR7ixPbDt8LXs6
gWjVj3mWPt/Q3il0woOG+0gABsxQTV3sJLXm/0OSG3cb9uJnpLOprq/qtqGkFvGSONqTVk3GVsR7
5znGNX3gBl/yLzwHqw+yuN/uYY8N+Ntuubl5wiOzGrjSLX40NFpTfd0rQbQpr5MlNK34hHpOVntH
wtiYrJI5AvYsIih1KrR73UL1Y3qDgEkveowuIlgDbgHiYWFuF1QmT6W52jRzu8AjTLR3jOIFAHF+
hSUCIt12PZwCRjEZjNq0TPS7D9ZacTvzawRTXMT1KriQ+YpTku3XHP4VWySwz1BtttaxbOabsp1I
yNWgm1mD7quMJa6BssrqYns3iuYsaMK1PUrlF1g25aH3jZfCyyscx0lo4q129OdF4WPhBP0mp8z3
0jEDyY1DvmDxRV7xC8hdQ/XBY2MOtqplDj7Oni+/VmHwfMenVZKf8UImq7/68kR8mLY8m1It3N9F
ds5lHsgDdL7hhpNhSXyvtrfoSMeteaCI0ikIgdEWBXBvGHOm4GH+wZmbp7VbrFUjtv0zp28L/9LI
Ps6KD6Pep6ezEU03nI4wTylOptEJdIdyaMDy9VQbDbkGU1wGxOsS9UZFd7Bf6AsvrW5DX/K6Dhh1
Ch5g/LOZ9+dT+4dO2+AjBD6NLO7k1JgNnwZ4cLXJDauGlepPeQ8O2IdloP6u4JutpBjlRbtQ4tq0
1S56z/dRv1BK10fXfN1/TmAAqoz/EeVUIip64pjfO9cDI5076+M4buKyKyDFaPtoHGxuLp3UmyTZ
OQKhXyU7Y+O3S3lCRdZH3kBx6KxlJi2CqlIkLKYhdRDz7oE9SU/w0MGLSH5HR6GTtQ4VbZryO1oX
/1/QU1YhcA8Y9qKp4Un3Mte020MGowl7CmrcEDwmjmRbQFk8PaC5Z6OsPZ4wBPSbau1GwvFWBMeS
diE04yz01VOyUmyjzIHFq70fwIc96pLQXyzapD8qvuzcOeLwd9cVk+qlriKaYre7F+rwj5e0h0Ga
iKrFy+wvLhrWVWuMedK1hqoL33MblYrhy2hUp14JxUXsaK+JuNvUl4ULLlS1SGG3xU6c9kIStT3g
N/J+UlkNWbHDlkMy34ziaVde12HfP3V/kvVW92O+L+zDrAuVGmy5B0WsZkiuGYwsmX6+19uPDgQ2
AzYBXEXAr2G9C2u+mCzBfKr/7rJvPNHjqP1U/Tz63QJizarvO+IYko6jCmqIGBQvhJ0C6ZaTESlC
nZYQc4qvuX6iLFpugkMKtFky0e1+onN13HfoUVe/Mhl5ylSA1k3mEzsqAEwDmtzdmh9TygqHV59u
KjN7mjdtPP4HD+9X6TiZwaEKzvlaErSF8PAY0sEiTITEVcLophap/v8yOTZvQRb4DXjyRVV63RKM
bi9Mcfe6+JOup/2Fz8FR2ZI7YZaQNtUm8b30S2Kguze42VT7usgbiZpCCuTJQgrLX7odkq+1Shnv
haA1llGFlIpBQRdmbnE4UpfYx6qYS0XBzBVHu1slPbJITRuufVz+o/MpSiEwaCmjvbWxypBq2twv
eFmUp8QqAFbuU0vcJ3Oszcxm/xByCigukfX0bsjfRbLWSBbwdiXefEX82Q5YeZOW7A7OJhuQqcPA
khfmWjE9h9hKI8sX10H+tcS9CKEtmAJDPu31SQ3nQXDW/75JZgWd0a3kedZsbh/MsE1j4GSlNUOR
5yFCC015H+LaiHN2jIp+YWv5MRAIu6VNCr7cTjCwVq7GhUnT1boDqFAmneIwIESkRsnpHhKJMvK5
6wtCWMH2EG8xrdX8jrbzS3UOtQD3y5gmCF/qRylp0PXPunwzCjAfJcHu0Hqg8+euVagXxNEOhspB
UpI0LGyCVStm02SmVhRytgXUfZ02oJndq/bul1hxodUtUQPapZ0TN6GlTdO/qZ3ner40oGRrrZmQ
BbAk+CBBPaay+ftLFmUJPO+c4pQJkV3gaUKjGgleHf3z+our/S3zHSDK1HaiLi7+dUabFAc+/qmW
iuDPTpDWy0Fgb8d9ACY+HC9K54cj3lNmLXBSpTfgUxLMOPcwsx85t5GsJmXLAPhVDnJPFy3/IrKm
9nx62ziN3vz7KYQnYb2UTxLzO41e9guw9XUVE60/DGhuwdBhoYcI5sjRuwG0VIQBakcOFrYtJxp7
JCKZhHcrGILI93OdulVlSeyCj7ORSfDbrrIitw/bozJ61dkIuk8Ru4m5ZnKsyR2Kk9HasC7g/f8I
82TwhqweK1vb9Bnv40bgz12qNtAZTX9jHi0RU1Yl1fD2pUVDOGczJ2UcW2q9Ej6ZNk1lEicHul4g
lpt8hq5V2nz5jNpPLQftQeW6Se88FBXJ2jSRZw558EUav9rwhUxkpKdakEBNUWYW7ifFp7wAbWCG
JEKBuicAjY27bW+O5XOOVp45i689ihsegJlWXhtmlbEVn08ZDGZekstwOE1xhqYrPgTbh80OHKk3
PAAORaJ0imXX4YycihxJL1/tOrxD9239b4brVhfERumMe/2tyLDa3o51Mux4svE0aWanUnkuH3xw
qgH84yOM0xVG8Dsx8pctGINpm6HnWD9/ih8Ajcd4EvBuvgNGAihxQfO1dyEgcC2+KpBVICwcj+1X
Rn9U/RNMJwg0aIS7S6UZxEIsgNILxaxm80xAAg1mKr48DHsHv+7qm/A5bhlQzELv+Shke+VoETiV
pG3IcCR/9Jg/6xYCCK/ScLaTV6DDGcZh0DrXecNnyegZVfAFlaTZGI0BX7lOFHeoU0moL2hggNs2
ywcbc/iFfXckmBCr6koQZ5rNSZoHAY1311u01IZ9qpzQaKLfABLxqOGsGL/FoaREahlJBnDiu9w+
LFB1lvGtP0oAnxmYhQ0K3MzQK4089A6l3YZyc4SrNO570DbaFvOy1ogRim4SGpVk0N621pyozPfC
d/96vRszQh2P9IqEslwB3cjkYudFBwlKuLnFlB4UmS9kUtnMqAfAmJr+p1HmI7pDaZEey4/TSiwR
ezeqdHa+AvWfQaM2j+C3cFnqZz5DEUvPxXgL+uOhkNWPH6+aMmp3TCIVmDj2l/857N4PtwHI1/68
aJtXNZwzGpzsrwgqu6fkumf8/L72Z8TfEBQsly3Oyx7XnU5FdY4a2W27nghrlBD7nujmclzJgUE9
2WpVecsEFuOfVknqcx1xsT59ur4w/zKz48YH6i/PJj4YhPgpdk9tf+0tHk90iN3rphvJ95tX6T1h
uXq0gp/9wEudwWOk4JJJqGR1mNCGUVvzMNsW4k78MpB5kaiKTflEmumnoWNMQiG/UfCIiTSXboS5
fxTNzbrOTLJlaMIZxqFy0dW+msCx8a3CVyTQNQQ4QPjfJPvNM0ckIxJgJ9oSDMEdtHubwKq+KbZz
mB+KcjmA0lY2xhBF45CBPYvgt2fKzyuu3PB+3nPKpq70qyy9dAsimvvzot9/i2FXXfgz5vOE2v8I
cf7hwYC63FVHU0qDxB1Wl+lDIF3eEbpkCV+JkBGhJEq6s0hycIt+dKAPCOTHlJrYLy6vfnUo52I4
PlCj47pfJWrO1kaJtB4sCjANeNlDInd6icl2T2Fk4HzaYBP91A499g83DQmlwxgs2Usx2MfNUGbr
0VrTGu/Yue7/TMmKQ0HkySXIqBRwE6ogxoUQryDnc+U1CkGsXpMaUVhk+f8a+25+3CKgi28ENoD5
Xn+I3dznjka98J5EV6a8vx+GB/oO2klS0CdsxT0aF//tmUfEUIybGtBJo5lznhlmXOmDoF+plTsD
cEwVh4Rr5qnTyhBwEF0NaWm94rshlgjspbdEdWCF6CjzeAVdl93BKXmFOunG3cgrBkCh7mDk4T9t
nPbGjxznQIdfA6+W87uqf77C/EJTOqAPV8JeTFjEHDyHa4ABi0Gy6drSX2TIkmN6+09m92Nk2/na
7zdQWfxvHHP4woOcTVCBO3Pb1w+LgES4yXx55EuYU//VHfLeTAA1/yAATAylRE2u8M0meOB9oPUm
jId15UC8NT4igiq00QOo8SS2O4eHI4UMauLc+azViLDJbkoOT7wr0BYBCI3SzP/FHPJa/dQTYI6L
U3R6EmQO3kCqKpFrrQ8OkVBKuT8UFmgbp/lG8iBeO2JmgzZCfUUONw8ffEfkKn8doPDja1UERtos
jZd98Mhi3qDHshL6bIfmRo0mfaWel4bzYPgBbBy6LsjJGd+1ivehm3+mtK0GKP+o8QVvdA/csijn
CXNnTBlAqRJjTP2fF9o3wWi7orelo7x95vNlLa1Na1jHCGPTZTjIIIWZMYe4K4tswxGShVACt6bq
SvhZDfoxq3p0xwatHz2/6PV40OwBtadzItQ/b2cg9Ejsz7H6f2NHbGA71tH6Sl7LawxiIfMDCWvd
CXn2NoeVUWLV+PsaYJRvI/yULqqwtiZqNgkEOI8X4HEL9viN5Ug1XRj+hN+BrFbEwGcEKCUEiK8k
z/AAwsoh1UfSF4q7XVpLsgqB2m10l5gri+4mxvFw137TWTL9p0K2ndrsKxzQwPxs1z8LZdfrw0/Y
0wIGfWkpEAZAqwG+XZHMHWeSW8xw+lus2+bu2cTgb4iUMtPDZXtyPbegiw3VSkrz4b6XRApHrdbw
lP4oUZNjY/nJ4Ut9033APWzWm8xNVELkb1a8CFMpwxHugWZpqRhYutTqTfeaCLVAbqosYydwH4Of
Dg23rz6M7lV/K+MZEphPMgcnaOd3W4zbnhM6qc0I86ALYaT+wFIptxGRwCUHcJ8mQWDCAqAfe8kC
oyj043Lb5hoVcjfu2ZPF2W+/alYCktO/Cx/6fdh2T1PJp6ZlcMQr3Z/tlZPuyw091mgPZEfb3ySl
vSgXqT1pMjc6WP/BOnBEpEjv/81DuDdEmwmF7GeOPLgNqKqd1XGxpNhcZW0IxyGt+eEVBhvi392G
41yKcSo6O2DXr0rzh044iQrd6FnBaf133ZmZRbVUhGdZqk862rIJdXsgzqbMK4qZTePuG1nCRHXB
kTJEDY5pui9wWYCEDt4wJqoC6HYFOob0n29lltNvu1Nz58UrGoEqEapeAiatWFcn9ECSejwUcz+4
PyVd7r+z7xFQ2MUMuajrnPChq/JhHE+tYYaiBWWOOAqyabkyDEBKbrHmstlapWkC/C8PosR2DcKE
tJcpIs4zYbYpau+dax4X/aKUrPRjxWT3zBEoY08ZbL8W0kBoIK4UUYjVeQcsg28l0zpfwYpZVlTo
Qb2riPNiPDuroVvB9A6dJTzS2VfcJJJN9TAPIv6RT6TLu72toET2DJsLL3PGGTfrFYtI7oehwYKL
KZBHeRGVGTxxSaFHUd5t6yHcavU2B1wXUc7RyhhpdQa0nsJqmhqHmDU9vDG9gcWozR8ukzCgtkdB
w4BedN8ge+wn1Sx6LG1fBubKQk8H501u4TsINGTXZpF+3zsxB+SLrDlnsw0YcOvc2tAF/8200hvq
uQQnRiwwWe7RgxOX36+Al9TkSe0Pdt4QIb1Ktk5x3fvga32xI9LT76UZaqGHyj7I6+OHpIBCUzwy
150wcJGi6+BMOc6sQI7/bxiw3wcygKiHtPqZlWatORSGnSXasiFdQWGkV2/JBO+EbNgiXjgtTaAH
uDNxkenWuxEI8EoEAnwMjnbA0NZRuJvN7/2PLvmB/0r8jnHGutK/KzuN1OSRKe5Jcf0a3ZuwgVqf
DMCYEqqEinqCp+id3X082sEgf8+fELBqiCJUm0BTVG4dOnYr0CfwvXP6Dwvo8AJI89pA3aYMt87v
ke5Wj8LkNjyan2Es3fl7C9+XMllorRQfqUxu00LY3JffTM5EYloFugMfGDQoacaqq3XWgQb5xdfT
gxPvPaBshzG+7mP+5SHgVsL5pbcj/JBwa8AwT9WFC+YatjAD2gUygDlUWTF1GA8p2OTt5dswOozk
lkbf0mN0OZ6vnmqIgVi+FEOwked+ke0+Kug+Iw05XZYeO5eAlPfNkDq+MUGQVzIUFtIidcjnniHd
7O1Kx+9DvG7JjVXJzOC7uU//FdXdM6Vs+ceD24CXGOspkAD4OPFiwvOlpKEcxzdAMv0UKBkSuA/e
XVj5IrU4YLKgrm/q7I0lY28MK1FSbqRRXCMpmQCY3S8XRqqJlW7MtN1Bv2X3BLBOQy2s7p9cMRmz
zX7AblVxJWNC8Sw8VI73O8+faZFgvRW/8FAxzuvV/nPKt+tBNT3l00xHcNwWIBFA5ZRiYCw0CwP0
jKCDOodyw6bRWZkYp41LTzjHTdJjj4xCuy6UjTmUbaC1S1ERc3gcz85aESLK85aa4xrXJEoJHmUD
XVxdpJjRci+ZK4gIRJ1cl4kRQJgvhDoDqrvT32qdy6H3RoI6DtlQYlgqKPv+vBwWZ/kRGpq791XR
H426UMqX1oYrsrdkaPYkO/rojQpLvjfD0TLa+y6VEch1XqFXY37eiPFLJWh/a5Ou62JHM/L77uct
+qPrBHgQFbhvFI6/DPXyWSHpOFJZ0ZFePP9UFHpM19Ff56X4/MxrDjF5Oci+9AQotVFxuZBx0Ti+
6nFlj1bSyvJe0idDvh41SVZ7Z1fcYi3hBn4emeHalCRJ5a6kWmAo0EGDuIwuBc6ZVIHQEgdl79M6
ShoxY1UMWPf0HOhsbCQSmGr0LfK25S6App4vLgccqbD3cAZfnAtI0kcYTJN/dY1KNeeBZ9YU8aoj
mELZEHpy4PmRRACKjZvn6IuOlLZoNMncldqHbwe/9gersosunQmJFX3V1hGLeov2IPqItPQa3CkX
/xCgFYIX6qL9bdp9RKHkM+JmUmpF/Tu1ETpv4aqocN0bj+Vi3unVnUr/o+3Q35uvvRqN0s9CMLaY
nv8taGy5f466j0uQ7slGGnhyJFxC17ZjXQgNxrfJJKpcGCR2ZX1YR8+XYzuX/6Der3X76R4o7U+3
g4ZEx/p855VgPDjpkFcRZztIZPJz7oMrLhCIJN9XCYC/lN/zDdCy74n6srYYN7KROnN99WqlWzEQ
8hEwG3Lkd6glpv6di1XuudWOQNRrsj7UA+SQd6ViiHbSDeYXGbbOXaUHh9D2z1KEC3y8By0zGBNx
OVPBYKZsb3/ojKaKkx6qsxrwyaxJdT2CB1bshzH6icV0jGWddyKJr8gFb7H+7qC59wemgf7SXb7I
rYkG4cD9rBy3TQfMAetirCD8f4VIjsGZUHZmKwrebAB1kXw6LGz5Cq2rvR0kL3y9QgKhbrO4U06c
fgI8krP+AZ1xtu07xZg7zqFms48hxYQcDR1Hu9qsUg7Gq7dGBuEXxoz3ZIvkn3oMS2WuNgH/XvIW
VzK+OX9nr4x+NUOiMGupmDhJD+Ry4wR5IFSkm7mI7EXMHPozE83vGfhw3YiB7gYN3kaSwIVVpfqg
yPBeMdeJJIKQcV8huMi1mkfK/cmgUJ5ZUWXR+Nb3PhMRehiDk145jnTLFVI+mGiEtZhOK6mOzy3t
4IsofK9HVfpPsnfdgwD1+Ji+AM26WW/fMEdjvGXzR3toLYSEXKMVJ2uarfEKOWfkRSyKHMG2y64L
agna/SFOjtJ24N4pSyXkLaZGAQkcvmkZqPSaHSGrs8hE0z5UG+6TY026+Sdrkd+m5SLpCa7501gu
b6iO9IBo7WwgWsC85OQ1Z5q8Bia5Pv1ccp4RGn5k/gbr8XG1sVi6fneoSjscMWjcsLayDI6UvZBu
FFI98xLOOSuZxotIKtOVqyi7T6xpPt7pUtJdPaqwWPQiIw3RAn3bOI14Wojn3rgPn4uSJr/Lo5QR
FBv6VXhC72ENoh2JGEsyb6lSwyL+g+ESvqGAG3/xyoq0lNMx7gqFJCq74TtBJTeTZdhUQLSoz1hC
RQ8FAOqxe+l+xIWUjGFjOEes8cBzNoALX5rBXB/Jjz5d2pUvRInAytmReKwLGoLQmGbbMQjsMhQW
g9OWMhqqfQ5r2c6qzmTeuwZju23OwPYvnCWO6RxZ4zfW4vupWy+TiAGYz07AgXZ+k3E3pgC2VfPZ
pl+PlTupiR6505m4bc2nIyDC45Pr99M2HdcOt9Li9gk+bLjmH3qyQaZ4mITzZsaKCt5PM7gdKm7h
QoHNfG1jzLroj6HNlnM+fshXKnqVIrY1UxLoxjjuSCp5D1K427KbIuBG6lpLJgC2DFRI8tqIwSdM
u9GW20NuVR2E9Z3iVZZ1oxnJldhXzNF4zoJo2RtiH/AhUFh2FgdGFsSrCxw21BPGwO6bcIzzdijv
MTuNESrXNGMaJZcbMeQBfhTRELl8yR/mTbnCiRwnTjrSZxEYroHb+1Z5SuGjX1CiGnjKXs08FNUU
4bf+8ZfCdY/8YyWTCptzA1y2Pg+1SJHtWE7JooC8FtSWATyY8lFtdxTZSfufA+kNpAjR5or5MUYn
G/QUEoz0qeyDzt7lG3PDJGtVHlLS8NT7nxPdv5l+kfejpttqRSmgWVmbhgHWXbddh1VuIkPGOP7C
qIUPLp+YKB2h3wSrWfKLWlmbK5NrPdfkhZd/XmSx/g2KzpokFMmCT/rJMjgay0knie3IK4FyB7Y5
yEal/6DYACeRI6QidLIgnA/2qjdm16cabHCzHy9RyrezqM8vovuLMnHWTFMpxTCQlMPzuFdiGwks
wrzOjk8FlnUupriOzSUt3DpOvryqh4q1PGQ1b9NZ3n7YqwJBtxzsGn0rzOP9ojJ6VPA+dVzPKGIK
gIniD11SJK/poNgH7jyfzkhdZye5h/NfzAhBp3gTRbozFYsYiA2gXvBFZ2i5AxSwaCEcfrZ/WPWy
NT8ddbeYeYacPpuHrC5yWCJGB+p1rX6fwhDXgpf9DNQgMIlPiNAOjSOPwwMLC0VBalDx0ESEe+uF
e/1Barki7JGlRpWiLbwhs9aSdoNOBAd7M91hayKqRgFqNHETp34eko3D5PEnIsYOOwQgEFrytibE
0+tevfGHstg2F/HBIqM6LjA0+lfuUOd7kzg4zk3MR1BpEtUqFAc7PH639C+w796cnVBHzSJGHncU
Jt8/tCRzJogs/d9OAkLrIShgKimIH7YKkA6ayQZ8mncU5VGQ0bHrgUklXCn4kqrcy2LfrCLWsioH
4bv7n+3f5JbIFX0H+UrLhLZQMJ4KNF9rnfHiqjmTWtxPXYz0ROhYcBh6M4XYppDgkCt0wBsLNb5D
pNoCisNFgQy3+NAGj+MUyRXJ1FVdTNxiyKuovYuCJj7tN8iKb912KtjpwIONyOA+CQFOEfmYH3jS
eJB2br3i6ndJ7Tbtfm2kz51xVz0Y+hJLuBzYRiAxzO3HWGnewG2ZPU+mvWycpT2GPfqdeU3UNmIz
QQIwdYbiTk27Ncbc51OvkWVFfPju6OZ3XtwJFuD5LY+G2pjdYyMBLxaq+m8X9AIUZYgkBSIKtV4o
W5O4JQAJMlRbgALq9d1v+5WlNVGuynInm4X2wGFTdDWEiNE8WvLkqddIb8e+03orE4C3lsftde2n
KPtEEa/IEOtS3KdVmCcDokFk/L6EZym+b0v7kf946pghORzrObJotIRYQPXAaB322IiajWT6lBfy
N7BUOjFDAqdGVroafpA8VPPDmmOleElG6WvU3DB6f3ZEt+NzuYFqPSEc79/d5o8/2SZ8IYa50JP9
48V4UzgczmnSLv14WqcoKHJ4HomrHIKWnVtVBAyEl2OTRppPoG7/4CqqS6G+pZneGsuRS8V/qzT1
QBwdGrpso8LP6iFoY/bVGpIi45+UaXjmfmPrhS3qBmIpjYBBlO1NbE+dzZ8EUa9nKWcsPGap5hWO
/xLcyOpWahEWo+sYEOMv5j5kRt/O+6MnBcKVoBZ+8XohJiGcQzfdQ6gEK4mjs6GSdpvh02O6q/co
qqSJSc2+/tNEBjA0m9I25xHMcZKlwaGVhqK89G5BzXQvRPEHHe2/bW6zKqx55c/e19LVGCfbGskP
isK+8wE97SJXCOuHkRmnLm8f0d3jXO3zMDi1RD7a+BzFLRhY/pEkQK8Z+u4AvtYh44XI4FXqRDe9
cXZyVPif98JUhG9H/otbcgLliFsgc14ba709yDVFBu1jiB3SC/wbdeRUvAjCc5tt4R1SoQn6FvoV
CRDV9ZwX0HEaODSplYx42AeOhVr3/UsWrs86hV+T4egN8qYa+AFLRFTo4fISo0IaVe4RZVd+N1fm
PXkWuV4yG8xrldVnx8z25yAh0s2xJh9ImunYQc3KdU1xFdObMZgXxLd1zXpCz7WLpO9OcBaBZQZs
8mPH0JhJNDIdhGj+gucp9KiJweBbZukDwS30TofIiT2ly7EXQjUWhQfMhrmTjFLqAbpojZ/6/T7G
pyA2rzO0J9FlxtqxYx1I2pMofrabq33Mp6ZYpqQSrN1y05UFBOhEvf7eeMZMZ1WVw+RCV+7DXaI9
oVkrFvM2+Bv7r84aU2f2xM0f95R+rTLgYxYbfI1lUsNQ4lexlveyzhW2eynVtAtnIDZa4BhwLI5c
yCnyh8sw61hE/x6n/5fh9Qvbi/IyHJbwvZXf15rEmu2nFz3ojMPfwGXccj30l3TzbbnE8/abg6VL
prMe28lf2K+2Nwt6OXaxTEM5ppULM7KTJNnFXwaSBG9Xs1R49lG0qe6NUPerpnstVMno2iMCpyT4
FcmYp6TWxtFoJmX8tU10XqxzoYlBXg5V8q9PPfEw4CNsAq1ROdDLFkaJyP3MJP5ornv85u3jXMiR
RWVIf/dkTa2ks2FsbGvlHzzchNqNGO9D/GMhWbs/Hmg7CskzkYDnKVZJkHFkifvtCzfLVpCq2bjR
JnbxTo/3tmwgoK5N2usSUnQTLfCyngm4WM8M58txxkh1X3vh6GMvNukv3UtgoCs1wRRfqSNAVpvo
oDDt61iH5acw/S2u0Q2kfvkPtBB3bgfHw/9xDRmqEJezf8jxsL5oii6eOb8bcjjWZnqPSRT5GPIX
Yg2AHdgQZzBcvIq9wOxfO9sifyK04/KURwC24UZoG9erUoBLL7Ca0D9DOck6gRhWY6RFtUHOpdR6
Q0FVtM46+T6QTSuDlccCfq5k/D+XAlp4qFXlG4TfE6GRC/9kuZXcjt3ZPmU+X7eYlvplDbCz7gwu
Wl2ewx8W3yLYpO2rQeAp0q/uuifJxUXVUchqhDRz/iCZM+NdjIjWH46F41Xi6dGSchP7EfwhzVmb
YYLP+F0CgR8Rvh7vZvkg4nc+/5zDEUNkxqiKVjhGA5ANnraxXzXfk3DwKAmyNt4s8LPcyrJeuRBK
/GoUAxUfZh0Dwv1/wOEC2XQ+SlEzGIyMjqI8Roo5XkI2VhINXdLt87wKnWTzvFgoIz4Hw5BZjT0J
r5OhWqCAXjSiTLhHyPZwY7rf0WHzVNgU+wHzrBzy/3uLCFKs4o7gacRLtWeFhK1as4VKYhUjP8GR
aX4BJKmNPbvy0P/1bfO+31l57W61WPkWffAQ0U8zjnhcEAJP+2K7tBJyPSw0TwO4hbiRuU/QkDUu
6iQblqUl+xuJAGxj5koxciv+zISxzcmKQPtrjHLJCC2aY83DN1MV4r8qcPrSuhc7pbJ4T8i+nQsc
BgfWnd00ZNlzsQ566Pw1BkPY3iwvU3kVs4cJnMxMvoJHBcrQ4oMVFvlTAQorCT6XSw/xxPAAMCb/
IOira1k4ljBm67eaYRRClpqjLQ1FQ+BylXQNzqJ3FbV5RjR/nLLZDVtngtPhLwiKOh8H2PHUpIWB
NbxwIWckZC3jxGwekiEOwaMyX7iFTn0BwvPlel9j25grVLRVB3vhC7m3e9Lkl46A4Mf6jpOcyebC
d9QoqnqrdYO475nA/sC2HpOkZkkv2YvxOhHSbxqS+ubQ5nDswG7cyTwERauSHRd85E8viSk1fL8e
jK+BlJm/Fh9fINtEFKJ6IutstwmSh/gHuwMm4BBLo609UU+Dk5wlhQp49gRm8AST10gm7QjR4RU9
eTmzX3LRefOchRzu/9g4VplDZHLRbW9y3UdKdAEgUUyqyCoot2F5nNoE0DGLPm1ZlwF4d5WI+L3+
ctTUT6SOaGd2QBhMB1iDvXK6usL1NwTTtEukP/S74KXS//edrhv4yGXQrU4IwErQtGT2Su17e9dD
qqxJaS/MrtZB6pItokw3AQcGzMG7gf+Yq6jMPkPJyxqfDmL/4EaRf3U0c9voV8tNvCt6+aQZhkIW
EVa06jMwdxNamRluc78Qywau1BEG4fdF5QAUgRNeq392956C5N3sR5D84037QfDBr62j/Or69U4F
6kSKysgfJLbVrrApNlT5AUKohqJG19QG7waHErn98p0oCq63PtN74hQWIHY7Gk3CHGeut3mjGZE+
QeQq6/jUxvyEFrAa/cR9rGTDSeNaGhZGlvDNS2kPiY7fA8HwuHT7uk0pn0rHFTwlgXY71eO/ieUL
aBs/1EWviNKneRMnpIPWvGbESEdbrLn0zEa0BjX96waKnfjMcYZEv+JkoQXnMn6zjaldhiX6yF1i
kqLKLr9yUPYNQR6MylW+2DuekRGVTx2uOflcIlFXtxXHxc+bEBKcDKeOUy83jLYat5rl9ooewvdQ
4lewX8cigvP2G9Uq0nnoFePTcelZc84GH3/P8/PU9oh1F9+TbX0MsbAzeXAFEqNCwyqWBbiwzMQn
GYGm39qSRw1tMWa7OIyusOI2rtrDX7z76fS9XPbiDdKdO4Oty/YQK+cQY3tkE+y1Xql6EKDmI360
OZ5gLA2E9Itdz9Aqi2oGQtFDAne7TqfaWRxKs1whWclh+Lg+jAxvqYG9CPdeuOSOUkCIG6doTaQN
yEIjrkOSJ1WUhwpWYSqoYMKw4h6zp6xzSwni7UIKz+hebm3mr9QKZDuEN16V9c66lQBuwsUUonrb
MVODv4TBjzUBzy6y4ubfNElsj6yeDPkXGtRWWpn/udvEW4UR23eG1/JSlAGe434KfD1Qe2vFO1JI
1f1JIueaL0H1bkmIdzPM70LpzDJ069Dp3fFgGpWMY0mevi9Cw//nl1tdzHJ2FaneKCKcEx/++RFK
oS7At4zK5gdgMQTFVeFHkz+JFyU0LVkEARl0d8MykZhmWgYTkSQzSIPXavfJ3//+gCDsAOFLeHd6
V8+KMvNqSIKoWkXBwctfLbf+Wu8nfSAK6ioQe0lxWq6AZoAVp55Avxfl4AwJFVSU7NtJqYEJLLHR
YPzKMY1sNSllOEPzYe6digw9rQPw+MuJ8oOvq7LO2cJpCEC1Y7eT/BSRdV0J+mZ+SphBtRRDFWb3
f1FF7Z9ibLALns8hRLSoU6+HFTN3vGkaJDnNfrE3dvBCH8hrGcFMHOJl6h6sWImeQyuAeWwdTubC
C86Gn0bqUQeHZdc0MBPxElvVxsDrySFojJfr05itjS9dNth/+eokBHQpVJYGckLWx8IR7K+Tpdve
9/SWdRY90CXP3bLdPIN4Fvksr9sMqoqbJpdHeYKWb17wl4L171PtDMRR/E9bImv/ofL8l7DhPpVi
NSAavlH5gzJGJoQlL3TeeQIPAK81KzVTgioDI9UGHUTY0ON2vEz0LlHytNU6G3Y50zErWR+ubuFX
C0OfOMNa5OWVdKjsCvhjSpgRFtIF3GYetE/KvhsRSmcPByPJ5qzXzvLurd+JLsOUn8/fztlc8EFE
ssRYnItjPBS/HEUr/Cm2NKkKetNOrWjfBAwEqhWonrk8/zGVo3Lhs7m7XtALB0ZJCvQaF0BWFUIj
PtF7JJFy7GbiIdhbeKKO48jXUdEbcU5tN9wMjrFKj347OHD3sx5LEy80BEPMzCCO10td1/Nq6I1r
LwnO/yqEoTrPooySrTNIaVzacIe/h1KOzsX4mH/IAn3K0lpcoJ579boBfEyASJ1JkLRxz708EJnN
fNX5JTiF4DoXIgJ0cjUxxejYVg7C5rD00KHPPQ8eU4u7O3G3VUphofWxGbTJSSRg04bM2CCjjNwV
8VkJFgPEowSJVTf7iCKz0SbGlu8zxjNSlKOudIz244QH86EfdIda9EFXYs3+WIszsb99lnzqIFoW
NH1AUhb9d6rTAQHsZ8Pu7goReQHfs+5J/5sxsLPgQ+ZJP/g4aAgiMmQipwH95vUVRuOnKzICqCPf
RR8d7qYQ3n1llsNxcd2JkE3FACBci1pp8dFDzZaqpCk3GkIkkDNWgsGclQtMtRssdpHGVQDZ8IyN
LhCYtmn/VlM0BJbSpMRoKldD2PL6fJM7y2HbjhmWoDVuqEbFXQ+B9LmgaM9s3CeByFMqSensRQRZ
6Je/Awe7gxnjQudT/4c4z62HOIGVPt7HZDc0qFJX/xYh/nBfvXEZH4lLrAGswVUv955Wax9vD3wQ
l7eTFhGIkpD4W8iePqCmp8FekSJ+u1eKpPPJO+zT2b3XkitPaorNJ52SfQxnNdVAK9S1N7k+QbdP
uM1OMeFjnU9ETxgevf3dDd3MTRf+owH+OT6O0Izc4d7/OlVWdXZC2m6aoJsLLwKYCInS7apJtHXx
e+ym56W8QNyWj/B6VUyGtb+MmLwtBbeCopbUXWagbU9yUgZnmOp2XO6W6FhZkTASDj4+/RIgZ6li
n+2+bEJBJiY8ngzbisG+PGL4cZvbdsNWIN8EwMeTPb2M8tI0UfWmb1rM3K1tGd8zCz03H49OjFPe
onhaOb4Logcx8nY6Z+0KikEUapaWOrk32EYI22uE181Be4itVqZOCnkC/FLLxapbzhxSlsdkjvn3
xjzfCb2Lq4pU1tRj6+2Q0kzBYLv4+g+14UJ4PJM1jfV/aNk9j5OILUD8wImCOVb4Fd6kN2vQRadx
wWmy6ydQQ5AcKPlklSRqVYqbEVsXTb5R46JVlfL8OxKJZh20zwLOMPFsbxUgnh/5exrKosuCiadN
gjziHlPnL/4HDPJc8drtaiccZRhqg/fDJ263OD8HfgZ73lqyxZq5zlxyTB2Ax7q3feR+hubRmynp
4MLfyCaJ/bc4YsWf5WtY6tkMLNpyFnlKJz7sNzknc+WmGTc2Xrd56eSdayWiRQTGxxHLdwRw6jTj
+O18qee6i1u0baCovZ6CfuR2nktZdXhE5/CZJmpMUYBYvaL6wCn96aTX5EjgJPDC/eCpAZU6QuGB
f9keoG4djjLhkKudkfhqBRRAlLiTyLEZ3BtYV/YYvIe++IEwXsstbhSrumWElQQnlqXGl4hwQ/YC
aIgTQCsCFPtdCBYpU92HFKRvmYHsP+xmA8EFz7xwmaqgZaklSPwvRHlesMRU76LHz8BOiyisImov
+yGqP8FhA/Nw8DprVA6zRDadVYPwhLIaLdnRsjgd6/WEsUauRAkdK8Ctgp3eZlPxhfx3HwJspiaK
fh0d1twA4Z4hi3ewarU+kuY551+em1D3cpubJQowBp/VE/H8tAJnEMqFNbVCALngzP891NcoX1bo
fZBYHfGomS5Y/vLL2LEbImT5GwP6YWISBsrLdDunfZBFa8+oYnwPtce3pZk+AmjKKffuIDPhkRO3
QiU8LjixEEbSCepo9mSWSEnMQC5PQmnXK6D4HAJ1d8+0vJyqf5EewObVcgrhH8dqCLg30l+Y8UUO
lW6hSDUYRVUB/B8XOS2vEcF/cv++qmjphMRagHSGQ1ozyQ71ViJQVQtb+s2IucE2Rm8s4sXg/ASu
LmhGTM01OSfIRwbsjwTIl9AgHky4XfOIeeh6G//gy2KGm8LpdmelUPCZ6gF1DM4Sa/SJbTMCCRut
Di4ek/0wQQayj++4nIUKbKGPaYYMi/uG/SQl48J0b0uctCEKpwVeO6yJ6ZMCrvWzzPVfPNDAEoIs
8OxHcyW3S3mm8iK1Gz0J7oqb/Ch5DuSikQ3HI5pDmvlleWl0jGmMKcerB8935xrkckUnBF8z9Dhf
2g/2mealEFXnHfJO11dNpemJ6Lc1Q2ch73bupqnW4fSuyCoFCVHeP/nAHlij7VQI8ZWpHTHU6y8i
LI09zFoeO7cPTdyDlsM7QA9t9F5m8TVEgXyrUiqrBLx/XBMz0Qbe9Rv8A6QQg7xNZ4CO5Rw3ZXOu
QeECSvRjgxSojmy7dc4KQylm5zLALOTH4qQhTebdRLJQRsFzctq6ZKkUUpuUvknYQHk5IqdmMhLa
d4XJojpIO3t4oRmbjlJUAj7O4vcwmoL4PMlwE9bPa8ogrQmfP9IRmaHEqqwD9yDXwVGRntN7PwvE
hIqE4FnLh58IShYt1BawjaKgvfD6+/osuw2g3OeWvlmm4BCLKQyw8VWQA1E1FQGXbrPtu7eBD2QM
HG+SN1LrR2su+hVIQ0IHiTj+4iQF4TTEF3BLw3Em9MlSZQ8MFdgaQ4W6V91DgRt2LV1kcUd9GWvR
ceyDX7PWRRapJ5Gu8jq81tRoKAEt1iwKaLe4zSIgdMkAUY2HppXwHBSUFqsLP7sXVUrvQTr7Ldgy
2ue5gFbRhCjOn//J7RSaWGrDnXHM0ayWNnZYvDDv593c8v2zNeR7MEjnBehRiu+wJP9t9ZMTEdRq
7q5OpXNmvXHn0I4CA0tVU2srOmV4slKvAe1Bz2jfyW1KjwcrYqEnW4xjHK9P2P0fATMKgXM1T1hu
kVA870LRlgbd0o7zp3moBbmtNR+iGrLjbBFtJKrFXflkBLXSnTJebQmJFs7osDsruyW5g1C9A4Ku
IB2hOj4JCoic/wXPUsC2W2k/uf6OcD539UX1U0MtBfRIHEZ7ThG+VXRJ5mdA35vKrzi2TmWVswFw
p/jRQVONA13Z15CAkoXPTrg5zNE33NusqrZcH1gSx3s67oL9hfoKf+LcPZiVn1RzRHtgpj5EAJ84
jr/GwUySNBOu7j/hF038LfoAqbR02iAcCabP72Nz21F8umdMsLPLADFNPK9JU6CN4p46YbtxNpKI
u3r6EVKVstHvJjN52DXbv+/9ygaodJVrz6dUc3QlLskqNx0CRTRzSQ++VRizxfJ/s1rdeH76Z580
mvUK7LhYRuCFDlkzGODZ6OLZJzDeY7jS3uoanGwU4Gp4bah+P9oCmgicimEzIJLYcRZRDxk6rATS
e0D79U5qbNg1NSpcpiz9vmENszgjq6J9M/TkOAf+6YB3BdRNmxtdZC2yinHJPZ/GKI/kCaoaFfVE
CdPC57yNsv4wtj7pwra9mTaqKYk5+uTr5ZP7gCQjRpug2bJBVvgq2QyXUQgWdxKcdlH8VwV/d+L1
EhfZoG8MBiCc7rN4GkDlm7rIoKYqAUqkjeuH4LqiMammEaWiZhHFIe8a3RIk0GzwZfmvIxRs+/lv
w2Spjb6D1U53iJAwHdwgnqt6T8TUN08qPqn+KJoHXYibUAf/EoKhqEMO8VnUEf5UJ2uUZ0o/Xivr
hRKnaKbJ6Nn3BP/kVuzcvExL2mWKVn4r1XpFdg1jnoieXHHuic09GiBNsmevjNLWsMH+sQNQ5fY5
SiYGoSTgoHtfbIbiW5zv0QLaIrao6loo3j7xzZ41Kj4ffAo4A9hfT04T34xLSRcYOtmgCvfpNmNp
oq3STcc9FWNV9dm0KO2Pq3SyAO518YQ65tBoksGedhtA3csDoGXL+HBL81Dj0X9XAQuAwfzEr54i
gXYHQiIuEjQ16xL9+fJw0RTSPOeboeYgjOJ8cZJauyjOR/U2u7c7BhVfaIVbTOuzdCLoKkt/GhJX
7RUzOc5xWTwOBMCzDTga6ARbA2Pf7cWayUbBlduvgIyGgwOJPoyrIug7vaFtWcmqF8Yd21oa02hc
LxjPzMgP32g99NToEODzn+MGQcsDfJV8SIWfsGHHwV1Qaf/C7eIeMtHTVUdjR6flWUImYZsX6x1t
e1D8gZ8qKkFoAd/6QJ9NN9RoHgXDjIhK08M862gz7ioLPyAQeHYffdjXCW7jBr0qzkzGUOOFyHEm
/8iIuFxIVHdAsTweuFanpSXmFVIkU4/YiJLbCMALxDJBwEbGYiYLaUno3IaedGSGH4HgwTo2Pej2
908cmJYO+aArj1fGw3d2MDznnIGicSBJVWQlCkr49JozhBB+PPvLdCwQw0AZxcFhEynaPU9+y5Q8
4ug+zzz8A7v9vMnq02W3ttPi+id5+LoTvK864SzkniMCpcAJ01LnMrtwYZdRu0On0XOuk/O8kvBx
565qM6K6yU/xL9rbj5qPB5KONu94dyt5KNk6z6kWXM5IhVSbWJUJ+l+AcUqWOLqNo+iMee2aC3Vn
C09JxuJB8b2K2fMFKnbqID0Kx8/MBLc+BWyIQ0k9infl+1ldSbEwwQS+9LPkGBnLixfz2P5anhoo
TzRW94NymW9eRfM/GhzF5CLn4M2Ke4Up3oPblxc7lWk7aYIpeCl0JOAp+85QJczlaAukKUo2iYbP
7OmuU8s7zrsyV5WMvhiIYzXbMUQp1xxhYfpLe6WSunJtafZLOBlF0i6qBq8ewj+v8pCI9j9Z1fNP
4bmveQ0QpS+I5abPC67jRMQf3VDkmv65zjMFjsSYxVmshb1yRrMUT7axSuntq8sse8zLXE0wCX7K
DqoCc4vAA0CuKTjycgEDUDuK/cQMowVSiHQJYfVc24omoSP4lMZyxjZN9DW1TU/2EvwHHOGHtFHJ
y/cvNFPc+WU8d/Uc/tNKvc1VysJUZcFvB7JxEF9+7NSc2NUf90M8gf3RPjgVcm5rsO2JMrZg/ual
PnXRz4kp/sOPni0bQph5QKauMdbng4FV/7KzqrJECAzGekXFj8Cqvb0XFwqjaFdcIQyKZbjSYebA
TqsrSjBvhpYOBEXbyZxGRAQqd/SHxPrPDhStHry/wPVFbIyqpppnTq3O+V3qSSgPmx9XnaQBTGIU
ebAbLGAv1T8vDo7RXY/65Q8SYtMDK992cadRYL2NEXA7LFEYVuHh5i33DMohe+YtgPRAOXAAwW1w
7v/4vYXNNYEauSxbzLQEGnZYkYrhczFDiavmLjIwC6uZXTB8UviSIWbFndSsT7rMEFezTGqfrdhw
XyJmJAq/z0VSZkAW4r8S5EtRcbBGq5LpEZVlu7yEgypXTx/CFYFw/qSy/oanZf6G9jIG7xe/3Quu
N+upIvc6dVoH65CCy8vTgJA1pYlF6UUiOBk4tACOM7lEMgVz+RVkg1qB2rz3Cku4CvEzRBU/xYWH
IAkHuHQQFJjuEnFu/1x9bepJAW7bhSsSY9tO/mgUIN0YhEmNu6dChb1ofK/r5oaJAl0UReuxiRiJ
pXWwrH0MlhEQxLUggI3W/5mX4OoimWVlH7v7fzUE4JaHZiswz31Eumz9NQVV87MI6Eg8uAxvuMHb
l3Wcvh90G/WGBJIquwkvo/Z2CFAHPnT3E5Jx4whip53b1RREzEKBalcDptIlOsSF4RScvXv9J9bx
4CJXxZk4Ci6/dxlwg8XTLA1aIw+JQvMX6ou38EVkXAIpNCaGidOwjgt+KQyGHn9jR4hUPehJPziL
qzcCc+coSK+690X2uW9RUI0dGQsWdArxoOipCKUPhUxenzt8GK6J4d/TLAqbCRXSpE6D03CG8OxC
AmgyLzfnDyQ8ukqlJVkExZ6LBY4cC6uwwzdoOh3lwxfNMPxPyihpd3KBdWBZpJPn5htKzMhHl5Jw
z1UHtp8HVVTumPAjK6pGhhuVqrbi9uAdItmAVUrDzgnyYLz2ff361dQGTWEZ+RdMHLRAubPxrgli
hxLH1r/tBuAePUuXAEuVUT6eWx8sYTJDz2Y5fZrW2S4MqH7lvUZxGSldFbpj9+oMX62BC1s00NsS
7UGvFh7dfBtyGTqpUkNnEHKC5hBjYsiT/Ax8kF+SMr7SVgDvZ3627xOAxyXzI5brKyrDzmhua2Yi
9BVOqj4LFpIpVbNSUiErKzip6CwfYSF2vylNXD6wn/PTreKsY7GAdd7G7BTbs5Q4DkGTDLu0554V
F5UQsMsCt+Nxk9MrJphIwTkbWyEtMEggXfGl+godZFcByulViZ+Og35VroMffBGW8CRggaGR2eXc
gnAYT1sSO73nALwG+ZLJI0gA3J3hIHkx1wSOf/z3/utzH/IBphWU0gfGX4IaQwIBlXfYu0eaOjQe
ozot3QI8pEwAkldQDbVVgi+g89YzydoXRlqeVDOtTsitiRJKOlxVrSzAsVOsNWWmYhr/Tj8w0H2/
jPRarMTfGHk3t1oEj//csf22ab0J1chIPGMhY78J1GQyKDutAX8yBPIW5d7XhfSeB7pmsZXCyRyb
jSMvfcgVgQ6KCrNTglIFfysUdcrHcBWZ39xW5toSaabibYntM9XEyc/xP4OWvZ8Ko+Y4fdre4KQr
vDZczsr2yCRJTUoyeAOGHARQQ78tk3eoapDESU+kI4yFRoFcUqA0AdlmICTI/S0UZqiMIsRDddFW
5oDMc9PZmGg0act8NpLvIKjVMjO3JjCoz2gnFUjQda7huRI7yvAXnkQRnpN0BXzy0ukO9CGoQM1A
D3Kj66wsRr7WMlnJhydOAWspG5v+4ybfTcAlLOBR/6DlBrBgXmDlYda6cTS77wTYeOX2svMqe8vd
dJevJES9mp8ZCkQJvKgqrnKtGNCaudsDefUFznsCWWHeVgIQNdgMOeVWk9uV8P0Qovvu6tdii/Fk
515M0omdERHvSf/3P5KbimlsZh0gP2/LMOhM+YHZZ4ikGCGouOSNZPVFqAs6QcY21APnkOxEulql
mbnAEvkwNSEwDr+R4o3XdsvDXKHCxPv48lf4bbHmuHsX6nKeJTOiEXljedgrisGNq1IVEJGtbPTZ
ssQ/bHWsGibxSgg1t0X4KuPW5ByOro9U06Wi98fITubQo+u4ZZilxV4klC8FNjdEDFq1x/M4hrka
OhNq+bfBWC6jk4SPHm7ONKU76XkaoUx0i1uS6UfViudPV+MKyW4r43ic59Yh5V9nThSoluVAxumC
cGWReekLjd7z/N/Pes+Nv41nB85CBdbzNwy15IDUTpKeB9xszIFj2VvBC6AvKwWEhGJoeQWZeOoI
OIOwdSK+xclJnSiktZ5+42FMkJ3O52pw2XB4e0M7U+aUAi2NYU9PFiaExriobIfkNQuMvSZYcoOp
2JUHNHASqs/MyiIOFBza6NXPEk+jhrsygRq+7+w3VyVUUx0kTzZ9LfMekDzG1lNntyGVwarnrACv
zU+J8BUZ9bhLxLnemJOc5rxNdOGXJXHEFWv3VjZThBKEllDj8BoGmyVpkvxUEwkkf7/DE5GpKlzI
G3/kXjI54NCYvzEnuIaThY1eOoU6uRYMtGqmOWDQDG19Z3N3yTcOLl3usjkdNrEREI6Ps9G/LQRw
RZozNJU7qvbWu8pk47+B0PXWq0qncYUBdOK/UoYPuZk1xiLc6+3nvslq705OI56ws8QYIZUwymvS
WWs2te6+T/eHGd1HccEtbW8tMWuKO7H8ZVjLh4s4atBdd6HvyD6FwycPKuqp2hSMEhmTmmIijACZ
OyfKDV1fdmPn6jYfRXPzgrgy/cJU1mc8T2LoNGe8pt8gE7FZPwFFyd/lQDzEyN4lPv5uNeMdVYlP
lQ/QGKb1OTXirgsPr1Cn+iIHu7dqLw2hvRNigMQhduRBj7tc7wZsDC1dyWE1+0yd31e+Zs6Gqnwj
+sahEe6hi9tG0D5kXFNvshs9CK7J2XXGWg6EJ7r0L0EHcvSw9v9ZIZecTtD/BNVFTe3vY6s07YP1
/uaBfqE2eDNuuSSi/H8+64XOB/EpY/vrvGhmGizfCE/b2ZmBDevhw+YjEBiPwzeYD+kNZk8kyEAP
LrVL1ypm+NDwy+ElH5tiY5fBUigw3h+YU+RwtQKUJ16p648HJOPmsrk3vafaZ0+C6FpebwDL8ZoX
M3s3K131gOe0aoAAljmo5qwuIrN4hni9NUashpASuP9rx/21YGX2d4qlQrTVk0kxD39NflNkETs8
3qKj6YDl32O+aEoeroi2KX8TujzdO0jhSOoX7jvOp7/43HmOt7bAAPIDBxExfyKTrXWuG9M/RPnQ
NYGHgSc+poY6ol20zayHPJNGSFV6rfwwR4RNG7OreZnwpI1DliI8GZDH4ns1Bs8C6IGV5pfhNX5b
QdaMVpZBXWHXOoDtZo7JjXfZgOJqPHSUkKDDKWyPbGWUWb4TfQdgmIgAADbJzIyUA7nr49Obm5Wy
f3D1lpaPJjseT2Z0ax0RSl7pHJhSJDV8i58UdskwrwPxFHaJRDRKg8NfpCBYtyz71+SmBBYvQKaI
CC2ZxAI70Oe/7Z0Mq4sxI/uy0jJXhcVKoyVUcJUKmepP47US7mxhf2NOuyP/M9Wm8gASPLV5t9pE
NToCSYJVjyan8zoqMz16JuEoELr8xyw7i/uJ4CjptHZIZw/pR+UU4gc+utoaxDBrYcoYLelOvdWF
3dMxb8aYumPtTa4+6UN5tkJNkGNW9+YUEcdiywp9nIl0XM2qtLPYDXh5JumOJuTJO5am0n4NcJ7F
o9SchyTvRGFgDrgUeR8svTHrO/fFFhyAcUdFn6MGuMLKaZPd2tNHvNlo/+dKDN0ADT8oc68sDY0C
u1E2caY0Wx5YzpDH7WIxFhDKCjfpqSWyjBz9FSzL/2A9WdC8qW6YvzseJlz+YLOKF746vINMVJTq
hBcOUUeThRlGoTUrNzbvas3LHdz0IJuy7pFhp+eyOqe9pHiH1xkJ5MtgdKzpHS1LBB09fkEA1xp+
E+ah0LuPx7obcg6zIDmTrbj6+tQ24VeLWUUpdDrOSyLfUCRDW3Ybbv/9xwChLBQ8MUkJ7m/5N+e4
NOH2dtoVVlxfH99YN6VP+UyNHmFmrebhJG4yPTq7g1DISzmi0q3Hp1G4h9BECcTvNd/nkg+XKVZC
lGrGUR0SLIUAuymou4xzVBTEAEk8Xd5yfzN6VdKZIV6zy4xDkvNE8b9asy/fZcwepKD+bEOKW7mR
/FGRZ+UblmfLuU4zx+vMaN6qdWfX/SI70B+zuAY5N700IaFHUK2Rbwk9L3lnwi45Ove/IK6u5sAD
LHvMVeFGgBmmilcnKMeJgDdn8DQjeQ8GOYID4+Fhqx6HJdahDKNRptsBzUQEvI5h5iqb5pG31YYC
G4gqs5/bljgse3Fm52zV5je8+pGEXZfK5VA564KMyN3CRpenYtmtlGrjg5wy5ok2NX9X1s2wnY+b
iDLGV66qfXXcn2hRUYuyQSeru2vW2/JOFk3DqX4tWCW7H6PFrJ2btTXNa1VKspBMCWg9aMDuYaLo
TxOPnYYCTgUj8wWvIszjw/55PuE/LCwSlREGePJmAv54/ArqRigO/Bc1djQ8+0AYHK/hVI0h3u4X
QtvT8sW8cSeeqSllOcy3CN58QeNUhomvJdJzL+N4DnbvI+986IW8P3ON999xHm0I/IfUciSPV9Tm
DVfjO9Hs/qx0TbrPim/2Xd32uX+EqKfaf2YMk3u8iu7FD3Rk4BJrAJi0o9iCkngNXuXOj2W1jqHr
PrHOCq4qhOww4L7G6IdOtOoFsanhlexfE5D7qf/mgpBQm9XI0Qj244+vMjgJcA8cGxUlRx8XKfi5
ytid1fsCEQmd8KkUZmPcop1PqqT4HdL6FQrOwL7VwVjSnvKql8b9MNtTNW2KAxHqvD7vqGCkbrvA
66SNdbo+qZIEmhNOwqA0Di1PwWquUBko8FjY+HGGJNKB9PgRvt6Co2MfKhdk3jVoPQ99O98qQXi+
MOOlGhjOGHGynyxo8mRu+ztReWwOS0iauSixmQoAfC4D6+Iit2Odwf3SfDRCMaaZSzdR8csaBKNk
Gry5wCgb1SHjXJWNkKLTGqQSHH8UX2/4oi/bAZJszXcUxYv8BCWHEgxBmiq4EQqyb7U1npa4Dh+T
LKMiVdowrH4maYxCDCGTfU7YC48u4OQiZ4S/SYHvII74woNLqT18UOb5OM26dGQk7+7uMM+xAkiD
RQ4vrf6jPiPxDqZjAwCF1wby3OFNust3pYWgdbK06KMFePMzL6VpGTbdBbeA9yxg0BYhxX4FnCAc
dXSzSyMl/4C/tzWIo5TCm/Vq8Qoe3mTJGIPKgSf3dBkRjrKZOBMohBWuIw3qMkYobJ58j+bi4hZX
P/8xMGx8IX+V4Ac2pTjb600eQfizPXQSEBvd2rLR7TZCmV3YMk51YUwmCo+Do1zn131JKS3pb3jx
IXvRBflUjLey6Z4HKjrw5RAnAvJyKwQVM2Yo921RFCtT7oUb7oMzpqwmXsZN3shi3VTFkHMAf5za
+iN6m6smRN2TBV0YZVPkT/aKFWpXaT/kYQxCaqogwcNqD15cCYgtn7uZUGWlXKlIXz9zXT02rDiq
CfH/GBI6O9yYjrIR1czuDLAHZb6u4DvZ6ySCnsweIjVNy23UPi3ZDaXRyuDs2vf5Q0C7Icr06SFi
J/HeUbOv7R+1OFiKpTnWzSh1JD0Xgm18HKLiKH4na1SsJxfGyjotlW+iUVe8XMq57RF/1c1fOimF
CQWY+sQU4en9QGs4fMTRwXWHRoRTmWLKWJikwbhnIg7Ri8l15QZoteRHEVP2jQVN7VOuUiicTHRn
T5JDCD+ScvD1iEuMV8i8m9GzsVFuQ4rQ/N1ySG4TvKo0TTVa1NfWsZ9qpNUyGWZd2MYppIYWUekq
Mkgi25m2WuCZk2lXuRCIscwb0+1vz67yVpX0kDH/BfhWa62aTQ6VHtFQgw4AYomWSyw/Leg1zz8/
4o9CaVkJajwgO6QajjLOEa0L1YQiYgd9RFM1qgJF1ob/Ip/iZmZjCH9ZabXhkZyTFN0lUBEFvYyl
YPvTa0JjzIdW4mkrDTOJTRjoAb6HnJGPGcxXwk0jDK04olyMdsOdqr/1zDYaZb6KVbLce3t9L1Rt
LSKL/DD5VueJSfAGQh422U9kczt0NXPovPGyzjzMK/duK5tLJb9sjOc/Qm7630ABDl0Hlj6v4XqY
SUuyXTB8WHDRz9HtftCBrd9AMD7RIZoG/CBC798XFARrfNXLGPl9jpCld48913/Ys02LNYB2DiBK
lp3bEfbLEj9hsu156Ih8gaIMJ276D4icWR04U4tlFDFtUBbs8+AwDtO6uKk/KzgaWxY0e7+hJLAD
pPyg29AXNmeMMG10gsWzinnNSkOSs/1ud4u2cBDZ2f43VZ8tU2Iy/rtSFiAPhxmVr6ks+R2m7BPV
i/1U2fKtK/yFMwZULVpZY4J1NZXSWjXyone1pW9QZ2d/HrTFMOb/vA7lY9GZxVt5N2RMpDTi69w+
SiuMkxkVA34t+ajSJuz7MepiePso96/uef6Ubm6hc7olL7kH+Uu2h8kHKuyYH4N+MsVr4J+n1OgN
//yD16Bk+I7EHTHLHXcr+ygXkje/zBhwYA9YGHhTcOLwp7fers3M8a0VWfBQ1tfeJYYoPXDz80Ho
AlbBsXUBqy1HNbNZcq9b30wneEsV3qdqrjfAfIZEWclv1MPKV3X5MzhbtRhGQtCW1PzfpsbaWumc
3O+9A2AObC33dSfCPjO09gCRnD8149V/JPty0rxeukshV4TL4CwhipvYGfOD8qFpkvfPDadFk3bT
knRVhdA2t5Gk8BJwbqWSgW30aVQpfeXj5+clboePmadc1o8aHHceTZIHsoPtMHPM+eyIr45/9rL2
fnWxJrgJYt4povdvcZhUYxW1ooojg7wHOA8tEBnpcUHKrU8iQWCKzbCGwZhcD2ysCFBqWAyJmPnb
UbmznF6dCfYQq2fZtdl1JcIvTcNJs7smJxGl2d5o2FP+aI8hAXKsU/wch8DcXHYch5P5GPP2AouY
wZl6L26/gzXRGlfnJZIy/zm959Sgh0+TDHpJ9jW/AW1OqvTdRSgU1ClDio/jAw7IJUfmmT2EXnhY
3Qmivrf7ASvlKcYKb1uVgt96nQwF8yw8te2HHYAn8peyj2o7oPNfH0VqW4kOo6cKhymEq/0Hj6Rx
TLwRSm+bo8BvSiDPmGzGZf9pQd7heOPU0FHI/PEAj2N76j/TuFXDDMgLKiMlq1oxhBZNLQiBrz/b
qbZDBLBxfbyIUGSWStoYSapbPUcQSwDmLEY0DQNnFMVMcv3tPHYpVxycr3Xo/wEx5OVZfq10mmoX
6bRWheMZoVEzJw7t2RH17K2E1LWhwfvL+ePm1VfPEIjn2ujrFcCNgjze+62AJj8RM7cJw/am88Dd
iYUsisfpC0vemt/LEBsNHzION7dXZ2HCb95+HdnwmRSF/PpGL57s7M8lj8TrrAKlpTtiYFdbqIMQ
cdQmwQMFTcGJ7PIo5abKKZ+b2fbV9DtugDGAxltC7A0CTuvWVzbJ/Xw4G9AzlYHEA1gXRvzcyj0N
gwm608KOs5odhQvsuQ2iCCBPIkSNcToX1dfx1ihVN+22CVQWd/nd/ns3agUuXMWcjZV9Ee3bVzTK
TIUnM87WSsOawBShzzG8V7X4STkX7j8Xq72n1geWOdfcBTQJk6UYmZrHSagYFOxFtTuu3+vxyAl7
oOTb5CYji7QjNGciyYIfwpSbuDL+59KTcQ7xSRH7ANBg5sbASxm1dKjlXZOaTCcFIRxA+iS/fOdW
EMkGoAVh+VZtWuYRTLH97PDZUenoNZGlffQHRsqNmuze3gAbjyj/znJS1/DwifxWI/6jdBhjELzN
LKaivYYNbRG6fMh/P280zFl2rr+1D8y9LW3DOvy/BUHKBa1EvatJZkIlHPlMpR6LC4vr0jU/1KTq
iQGlsYYlkzl9hdypyA8XP/Bk23rR97Y1Voar9o4DYGjqkq2T/BnXVyR3zpcd2t09D5FkVf1u+q78
SFdM7LHXioCBxbbUPUvDvAI10IBp91d8H3DTSuHCJDB6MvM8qHT/1tfdGl3dC4cJeaTAz/5ztiUn
zasabgdyQA809cVxrJz6aCjctGj5mb9WkLkdin1cjywrjmMCXtNK/a+25F0LF9PdUo1pNZTjhqif
xEVybPUuol5OB3vLBxGRiKQLwB2o/eWuSxi8hi+VWLgtQMIRp2IqrU8mWVbq1Ptnr+CgJhwP7l+j
g6cEURyCxIqm61hMxIWo1OtjKwyM2F5OcxV6JG3nYCT9kT5MAoxqWVzri082MqOZ00f02as9zLm/
Xl1badMZLWT94/ZdSq0wf2KaSnQp+cN13KfqR3GgoF0eolWjsticokz1eREIFv6aLxEaJjQorOM6
mGwk3/MSx1nZAyhERIjjRJDeBVYJEhF0sxkrHH5C/KlFK6ZTlxheAl8A28JJ9NorgCYafoUnh6+E
pJfAwEigRMZYOvNWeySCj8+Atykclhw4XJlpGF7mjTkXB3jKoxqQ5s/pwCu00+B3d50Gjp8LrbXv
UO9V4n3D6fu9yujYbgGA67E6+Yk6BuVEoq62hl+zMrsuopdO84HeTngafYK+nLcNlNxMYmpDYjOz
F3iZOG7YJzdILU8vmMkb4uUEmrjxdDQD/TP4l3H7l6FHQALSwiwTNq/SHze6XM0nhAyglxH63vjs
7gUiWOipiUhdJNBLf0jOZ7MNRRgsvCfznCZvJ5pCTRML8bHYV6ST+E06wjQrfKRFsWx1QFlsJjzY
1a2mrIxsjy3w9VYBh3yU+f7kTlaFLgBlrOrpzV5FJ4CXr6vlFwgOnXwB2BiOvCeZwnRlw4+zSyWP
gy0pOHHA6wSgGtj7+c9M5NgjMoFWyhXi7E0nZkDrr7IG4P+piFaPSG8GEaJIsDfqmdLNPNsjkGyG
OWjQz59TkV/+vpe/YyQBHNzbdwbg7ImqnoJ/QNXwYDY/xx9SmnrnsklVJiYYK0e9lRQtWGaa4+GU
6h7w6ANQElOGbOgncjrvaY+iyfsQ1OmXcTK6/QaglNoykwPTUH/D+Jh4H4fbgwsaDoHnwk2hblmm
7M4v4uYZcAItcAILbKXQjmhaDIMD9Q4b/R9ZQZlxGrWSfUeR5LcQRd5zRT1YCZfzmp8l2uBCnaoB
VyHOIf8UMnl6ZzKwJPsSSrQ8GsT6fzQh0pBt+GUUFmkRpLk9si7+/r5DbRKEq+fnMcA+34zjCJED
893LWQaZJtKZiR5N+RDYoFlGcs/WnK/dKuCBGNzBLnkmFc/5JUE4Bd+LnAvH0T/eK4PPSJl0d+47
3WMzSAEylOFGZhTH4fqEJkBku/e7sGQyVf2iMcP2hqkmKVbZhj3A5OQnVPIQ80bfJPkj1trHJ38k
nANpD80SRa6DRBRXsFMpCzaqRnlG0JPFiYSXs0Chtv0uBb6Xe8svcesuiUhmabq4HnXIEXAnZka1
FNHwgj5/BonW1Pe4pPduz7whczb5tEBqQQ9ZMm+nlJA/x+BBLNrZStlHJPqr/VzJmigDySAJ4AGp
xSOVBSzYag3TsU+wzB0km22Drh9ZBMUKFfmRcz+LfDVATGxhtbwSVtO6J2HKZgiKgGRcfg6wJlla
X/dTgW7O8KpKIhE5MFeiktkYeS0JM29lTNu4M2ab8L4LjnJmxu2W6d2jQ7oZOLK+vuY7K5Wlh6Nf
uNYyWmvBkvVZQhKqA4VCw6D0s4KbmdPRM9+Z0KcKtKqYuxneaRTip35iqKmd/VZgLz9A3m/75zFg
8e/NwhTRAnzENI2K0NfEOVVAURR0jEDOnjJFEwpNh5Qpu0RJ3Am2GdePctMAq6PLRjL5ZozLIR+4
R2nCrUW8wO1FcyT/0mMoz7K7G75NODoIj78O6onf3wVAqzRmbr8aO/uIK+YdJqiuTXU8DtggJgqw
nMWuXEZPvmh+4LCGxhMCWTZl2QN29zfCDpbRu4V3P/J8oC8RxLYtG4tp8IDGO2kEP2N3BFi/eoFI
4fjtWAi/cF2ck4PNmQFXz/yeSfrliVUcIHBXgEalYSEaa8TG/PQj6Tu6TerJI7YB0iKdFKaZxJLf
x3neosQcoggUVD81gVYSkbP2DbCu0l8VYN+l/pQir6+pNepvR2b9R242iU7fiOntIrhLVFJQSTwT
trtvgIU5G8smEnXuAmJPz0cI8hO3QF/kqPnULLlTh+slcaVJn4ALORnPgUxTEELbVLXaagRiy7jS
5jsoQxcVCKGj+E1BBsNJqX8zUFL6Lpv2tSYg9cCrdM5brpk1AVvEbE5/fBCUhVvI1Ar8ABDPrOXv
3j9crRAkFcxESLD4bIvdOEkpYNZe86/6hz98YhGRhi05o2yyKYrIOGq0uYCb2EZogW9QsEKNMY5b
Odwfzyr0mVd18j6Pdey86Gv+XidlX8bkAs5FbKCEgALi/lMc+S6jlCdqoALBlv/FJqliqbt/texa
0vfGVcHapThwXR++Wvw+peaBdSwC1tFpJF5orCaItLhDXDQybX4zjKcfz4CHKC4Dd1B/IKsl+6rd
U2pQIEjhlt5hZXz3S5t4YBiUt3YccmlxLI4n9YBexetQGDz6DhpKkeH5KUZsAP+BPgDvQEAjOcTF
/emwqjIDxEelrBz6gDlNs1AGzyIC/lI6b6K0Z3bJLwCAfTzqkwI+DXONe/KGjSMJ71450cOUlcG5
008RpRsMCHwgrELdUbgfNL8l7qZpWQeLLSDNcfe0KIMR2e0Jv7XtPNHihUVKCnwgL83OYajjBcMN
89tjTrUw3kfAzKmJpF4BhrDiQLhfZvBO10Ax4hrdS3hdeAEIPBdRQh4T5jfew5KMCQ3iSbhov0va
C7LHGzbKIUzcBt/KTCXDQVdP9FTO7jXE2mx97AxMStBQgSz42rAkDGq2FhokYixP5rn0s23d59CZ
McYK21WrgncT+43g/5xDSiI7ofLLvinz2gnRZkwLgeIAm9OKPu685JQHV+pT64pnvZLcQxtMVbqV
cnIVvQr7VLatGqmB8cixA1++vQF3ZKDZx4xIXHctHiNnYKatv9A14vQIhJy7LN3loon7USwWq4pZ
Utgav5IqXuCpCryVXND3/hbs2Sh88m1NrI3cn17HzSc9EGYg/aUV0lgzmr+OTsQUpXFJH9HurPAp
/LVF3JHxaPrro7OLJRr3STRvwHssRrEWwVP8WVIAIF/RIJ89HrBZ1m4WwIX7eUmYFsYstrf/26rh
Sog+m/Lg7+jBVJ/g48zNXEGtRzS0HerZo+cmolDkjD7IlWTJeQhJLMFk63lgqic+jDHQOMvyXffO
KPiwStfZ6zSTkmF/hJKEDrr+Yhxx6u42ZIgK3zteiz+Rtv3FFTm8Ga+bvJ7L8uUIhGF5iXqBXKOn
bE28FAYQhVGcjczlz/mV0bf3HyZhsRS7paFCNDzKnOKTsV50eAr55NgBRQK9CPgDHo/jpYS2wVaT
V4M0fdMW7a7hXHcK2uIhwl1tam4DJStYPkq6o+KdPxojIhOZnPBCEwFWb2klZaV3GsQ/zdAccJDZ
wTB4uJLXQoulqvPOEosXhhquXAfYBVJgwOV0upNXyFR5m9+30l1wqXOLBOajma09fmaqgsX9arF3
YyOYGCLbqAT/Ga/UdJaI/kAgCNxvJNCbPQ+CPMmTOLhXrvpusW4IW9zD2VfKioUqU1prHKDca4q9
uL/5IXWaD8kuQJB/IGQfdsCzmTNH3tk6PQBFBLqafxOd9mUWy9wZvYB7jgvlFp9AsJFbnyywwI+7
roRUs/m6hWYOTwUH0T/Wxv5nvB7NPt+4LicKlUeWrNZPQu5uVb6zYqAcXrD2Ajiq82iTWi1mXNzW
mbsK6W/BMOaBFt/WAzJiSqW1IOt1Zuo9BCubm96R/NQyB6jTFFSLJV7xykTdhWEAitm0Gfz4h/Np
mT22fNHTEzocxfsIU6mfebuzqoK182yQRDMR9wVmBgOzHNJ1knKfx1cn20smRBmCV81YXvDXf0kZ
RHpqxKkwI/JFoSE+Pp0fkOvN0stOJKlvnpE936rcsw4QZscdVvq6WQdVEKMtU1Z1DKykcp1OZNLo
hk52d5TAPc6RUvIfTOg4Xe48P+VR9Yw1iW9bTj/gztYoQZXbk6NMVm4uxKpU15iQ4Mus5gp/GA71
Sh3iXNUBDjpD/CCMVc/akRK5zpI6djRdDlyB0NelVY/oPPpUpruKYjl4AgJTUe0fJOLP/Zn/dSs7
yJfT4oU4lpmxZF+FKKoU9HEKJ/o7Ldc4jv3QRHeSTcDeJgsssXzngEeezjyATH96a6PeSkFT6QlI
RqlWZwSAra170Q+isSN2SYzPvTkG5yvwwMqeCx20sR0JRiMfRqL195cxsbY0QifTXh/WDlCZ4Xjv
WDXmwujK0UHIdRKpLuENmLstadyAYrB3Zyi5TssEPzxJ0NrsluUEFW6X9eZh+F2z51Qp9HtMLwP0
sxOTG9IXnMz7k8n4HGJEleLtn9mkYaCkXGAk5O+cXY9EG4+/7lerz31IW5Ist3hfbwnfxAgybBDa
VXGJQ9UcQdiKZRrHN2IvNMvM3JSt27RuAy8fPJo3vxw0Oz4+vCcjT94Os2i/hmGVcdDSKHtD74aU
4xFb3jcwAj8msf4KrdFmhQDO5mfdZ1iyC0S5OtZHLduEUSIIK540TiV/prbHPOCfbQodlaSCKBB9
25daMVGJat4Zff4blvoQqpzuFwNrNNxzDzPJZyNrVbOugpTCZ1Ofsg49rjOdl5qFxcdKhTLCxZl1
zTVuLNNfJ9pdkYPIZSld3ol640q5seU30Ui1Z9cGskbBxaR6GiS/S0bmu9iHeMJ8FMNX5rK3ovWC
Wgauq1WyQkleCg7d7vT1/BzpyoBJXHLkawAL+K7PwD/jwBQBIRLmVs7KrDAfefQGyJMCG53p6maA
N+kxWNUV8fKg/ort3oZ3rrLwPc0XcoLbALBN1iN5WDW4VK4ScMpMYp0DcbhHmsrxf3xcSYi8tQ9a
brhbHoqVquHvgMKTwBbWJ0LsEtBg2StX7K44aJVbtwQO7V4t1aoDry42i7mpNjqgvQ+y1TpRLk8y
jXSey3VEkbejf7x321AduT8KCYxFaCxK2IhbTXNekRgjbi85+KhO/kY55gycin1a1hYnrRRzYtLV
ZiOroRQsANbelJQOlm0fgYTXpt2al4jB1Pk+dn5pEEroWIWwblCnYc6CIHonLOSL+Ey5EFIHYU7S
XJO8VSI77gt8S+H+HmcKuOmBNHvO9OEOaFFAhbBdFdf0LENlsYsqVUk+ZdSClYS0FEFhDq/LktF+
jjI3lI2T8GfTu+n9MVsQkhNOhMtlRkcLwEhQd9q5f27lm5fQDARYX7d+QS6KFh86SR5RnKE58TMv
cBB98U7hJIh1OJ5DWZ7zEKhm4Xy14qzTQaN4gGYcYMxXCnOuAQTCr4NPdrGzSKGGOK2SDgrCYwf1
nuUrs+t36RBr6oGrDrEMYMjDwLAi7VZz2QAsjQDQ4AWEvHybAjELkOFRc69DYzzizS3HI5LdE7QC
kwYK+mavX67pApeXErnyyT3UY0SMoGFsHgXySubJomJJ/WOyk1n6ItM8RNq6xAtcBqopGOGZo/yH
10Bkm16op/mOjd3cT9mykHGbQgKyLXyPIRAx3JkxeBsm5guKzqlw+q0tlIa2iBNvqwOsbH58rPS2
YXa/U+8ht6mnCuCAB0QEyCUXVar2I+QAScSvxUSXujP9JvmnJpp5R2+Qgj+xE7P/V3o4ldBk+TCC
Z7g+RxXvC6KvYJ26aLwlo7vhf2LPsFva1d+hZ/xv4sSEpXMK1ZiWGU1L5HQSeQnEEdBggxagOmBC
H11mVsNRFdorHN+bjyt4q2WOT+trjkT+l8rXHkrsquM4FhKeuO5vTz+PZafJFu5UGZJOHFyZK5Xd
ZoF8/9UQQJjT7AU4uc/uvw0sfwKYlAjELGcrykdy4tTumy6+lqZ87xr/8z6+lGi29kUUNdpby+XP
CzGuO3Bd0mOvEbV9wMC6TO61WMmdR8rcxlNhVmb4vdK7J1g9kdMaRikumAFR3zEob3BUliZXlJVu
b+HtFUDs5pNAE5NYUGKyyF2yz3RRubXItRYV+qbKut/M1snGRn9OrmppKkpGFYnPCN/vOGm3Ns+s
wbtt0ZzXfv9z//WFZz4Nsrod09mEo9bsflLaoMArO5m8uggImkurcwap3KOB8Ty73O9Qq6zXO/5Y
Wk2ERfoyw7uGidKInJZAaG1gU09uo3dAqB3h/mnek1AMsjbm4kpJirvZp+fgjjQ0QnQwGMrWSzqE
ULsY89KknOudpiMgJfBpwFLTeJ0mNU0PgvU2sL1IWf0mOIU15Cq+uyRlsXvtJxOgxGEw59zbWyZf
AqhcDbufKcVxKXN/kOy7gX2HCYktHRfp92MDw2K+ythtfCr7916BsXB2QJSKlx3uufWPUOmRg5Y/
XSvSxBUVfyEjps/TKKks9iytlB01viTKIsBkgTrlPVtIlHxldqHnOXu9r0teOGXZEp8s6dQRsTiI
idesPBpCxJMAmiVlySFuJmDjbLxasN8dfq/KUCV/I2HUm7Ld7FZU+lfHjaL6PSNFxsLpgdkyNmJu
2AAxToiZGj4uRu6o2HqF2nBHogMqcZ3XX0SzxSu8bgTcPTykCZS0o/6DhUkNcP3UNs+627+hmsL9
nwpdQQkbk7v0tBjHUN3UQ7BI0C++MTtdBuGCGWBQIarmTH7tig6Wu3pzoZwOPxYZjqlb9AMIN8t5
7yf5jnd7StB9QP6ziizxOOah4QX5ZtQoJr7k/3BOY44hax3vhvi0dTIsQFqhXeqPh0ewn8pneub0
cs8jYfeLNYjlmv6AsNptLlRVcYVqXRCxc6GPYnn+nHo6UR98+LqXkUu6x4iDI3tjN0dyRd6dZQKC
72BNZ+v3wmNve+hnKXtaHH0hwBLsjcc+7KeX1X/Q6sPlMQU64pnkuwWXAfQ+OD0JkyX+1h6OY7uU
E09yiLhYgm4PQuh20sknAWEGALZxhlh5Acv2AgLUWMVX+R9EMQHA46Hi/QAZXIa7niaz0er5Zfrr
O2HssEABk8wWvyJXb9ayhP7O0iQ/bprCbkrIS+HcQ7SN6YyV7EORafWSIXxkZMVpTYkPHCvn9o5n
NqZ1vpVIp7LdkP6XSlOuSDn0gyZZuYICfnvYOBNBOPjMLJp6au+eYfoffJxMfnljPttpop3aCxsl
R1sGGKT3kJSW1WHzj6bxPemDqZHR2v3CEKaUTwg0ZlDw9Tng5kdj9PWZhEeXGk76Cs0eHvhJhmBj
okphVUU5oSgMjsMfoP06Ow0U/QZuf6KZ972LGWc8jJhhPsGLDHx0fF1cDxk4NTA3wc/Ir0YqSKHE
v11Hids7NUkc5JNR5uCiUGqUXd1auFxNI4dDibHKTm1qlFtqT1jMd2iNl0zg6O1kAv0YeHP6vEDa
wiJl9K/6Ir7BL00ffHYsPhdNu1anY0MyuERHSeFVWAHKtm5uMDSZDRE8ghurP4qkoguYhm7/RooC
H7Gql6pu10spjTDXe973h/6pJLFUNQuld/FIaPgEAsar66FLyvF4o5vz9cu6j+DxRpDRSXSd+upi
MDejRcrLzkgY4/xAU7zZlR8tXL/7uDS5iUn25Be3uxNhZdTxOWmUTwxqy9ULzKWRBmQ/r8Ak+xcY
6Y3W8/pq/2hSeQo+h9D8hd6CxNu9FrWp8LYGIrZuq1gYigO7i9hfiV2X81aF/mf1V3wS2vpRZzrs
1X2gOm0wOY2pNzDELGFo0+C3eJcCR3B8M0+XAJH3FMwCs2P4Rg/Ep2y2+0uQPr7I9X95+8y6xsSt
VyZm/S4JkkmVf3ZvUZDp2enkz2u2k74BJRt/wLLKWgre8YVOX2FZxozPUM/ZyxeI4Bn7aONFZPUU
I7QnwOHZvi15zh2+EbxvKVlVEzm1JPYloXze3l7EBFlwWDgIHWSXWogXhWqww7Sarxkdgr4iXxP+
yCx3KyPIjmRgvqG47a3mvDgyXuIoR/QkLCPvQBdjLqB5TEa6reQtt0w2aX57MO6vhUpoRmkM2LPr
KbzW+H8D4cY9LTvocDG0yxqzQEIHBZfAVuT5QEKTAbMNY7CR3H/tlHAVsqHGBLZ1nZYMKe44jiiW
eNoku4LRnXlftkctylhs724EDxKMMtBjQvczj9a4snqIx20BgJmqR6FbQvA8VKxG/YKPk/P6CfY7
LHYFno6ZN89EmbK/HjA8S6p3y9PY4xGiyNSoRYk0ceYYk1N5XquosGNRizv/WM1hjjtfqirfERgj
Oby6ZuwDcMwbmSHfLEaOSGXlo1D6rYJxKg96kKx6U5YGj+mTP5nqAmmNM43zAJX5hXRKVuJFg9vs
08nQveq/r3z/K/eskc8uC1nOjX/sOEaYrq4ck4m3iOtnUN30MSbvHoW/6MSLFjN0r6Ymf8fUmNkc
dxIqMeVYkMxssTwz16GGHZRXTIimWBBJAOZkYYLP/iNgcMV5f6wDAw7vYd+AZZdNGs87QLY0mYhJ
gGD5xcbOTnxu5ffSZ9r+qIgoWy0Bt/i9G3qLvcmZP5pJ2Ad4C46EqwHzo8hmBwi2Bb5lUPOQMs10
KBWa3TdzJDbZiaI8H1Mpuy6zoHWBebMhgMmPEdi7TCrIXhiNothDDkxn3S6BIIUTmazwIapGVdW0
4IA92OstlXAYJ4xjZwGwvDSmSSYXNj0GwrNE05DGy3eGWjtT0l6BsVhAndYZK2E/PWK2GR6GcKJx
iWuVbvu/OZAHAro/ht+paolreEXmNKStuP2ZORHeYZ08QFdy6+vrd5RGz8RS/fHQZPGByD4jp00Y
DHKtgvjfVatDiiXGNHRjrNbJzLfloQ8wvGdqnSST3dQogAgKO+GB5pIBFgpowjyqHe+NDl5gz6G6
n6KfP0CtPNGNKo0/ogjTAl+1nKkP/8YHM0g6Mz2eXmt5EioxWTdPSQrRovjiNd4BBfCuGRzrIQDs
D6x4wfTMuNEYEz42SuaRZIHpaddPgyuYZOpalr/6o4COjH+I8RUzXp5ZdH3mow3a7hnu9nfMa0kL
Y+oTFcyLcqqxf37Vpg3CLHyDKIGXcTxS+illnZKaSrGYTGpgymTHwQtNYySfZEVunNQ9X9od9N/4
eb2zsXqN0clBeilGCbn72MMwaDWbg8Ms8/BbXd+km8ajLvbGqUiBIrAhlc2vonR0HlXxkb40c4uz
jGBg/FLKkS9Fzc03/u2iit3OPQ77iSfCUcglwr4MzE9MC4+/CqZTNx7/yunAYUJSssogKUk7Rq3D
2kBAGEaVB29EJTtppiKBoUqnGoltAvN+E9WkHwJUvyeYW18Nki2wGfJKwldAl+ojI/WsR6OHJbUm
vyTpjo1yHQu/H0fOmBttDZEFxdjkIV5kT8JMFmigs9GU4sa10G95oJd2oYgrn+DzYgdxVI4cC2Fp
PLYQPAMp877CedGHvNEfPFwHYwsfhQFWkrlzEdlaFq6B/k4Sg8IZ5UVffubkFinqVq0s7hr5DYT4
yyhnN6j0kkXdR0fmnM9c8pamVikdydAb5PD8xGGHB8NPRndnouZI5ZJayYPPbvQdqAX39t2NLI+y
vriKLbDdOPXBctg/LSveJ2lnSTd+JgQ2cndWARWs7TEc4KK6u98Qsi681Yjh+qEwYTGEuTVIl3ub
pTZCZTupUoh9eVULiYlATPtltUa+egRrfntVIbemBBzh9JOvKo0owf1fxtc20wE8repFFMpKb2uV
M2foLICBdU8TjUZnmy9C4myLX8RwSDzniR2JO9KW7MwMDvG2M79Z534gw8RzQCa7p198+wrW9gKD
x+QtISoyOCk94WI+VUkg7TWDWITQz9RV2n6B323X1JuSPnfo+hJnycy0k+cMHCXyWy77isfCbeNT
Y7kQrhiOvzLmV3ontplFncWhxe7XmI5XwmMhhFe4TysII17KH/PJCcTwG/rRFv39xvPBaj8pxNer
RcXMNR6C8r+s56ueUqvM4p5ZdhF29fWNQGM7M1KvWmM+uY9PsTE+CbTF08MnrblH3j3UV0JqkAGh
D8VFAGF/0waeq7Kyaf9OKL+EUuNKrTCS5psH0lj94dm2hYcQYxxOfIk8ApXiqIomaM0o3b34kzTt
W5lk31bYrrvMblMekxMg54vybl6krdDEWk44Ue8DjDM/UCjDoTCDw8vP9vwP0D8xNlP4VhlpRnRm
UgeUwaYAGln9sDb0ecOp6yF7jgJNaA66MRwZ7W5IN8qnCxwYj+j/A+IhC0izLDX9HxKDcw3Wcxbw
gnYyT2GMgpA9wOiPUCs/mYdm8jxr7xrYh410zgtb9MlUkwXnqbC5FHxwkhgFvCgsFrOcQppVTK7z
uiQwFAbFApE4zVaZXt36ag62jks/qR4wtpKTMlBjYVYrLXPXiAvRJ2LwGnWNMgGbIJdNEkDS3ciM
aok4+8ZaFk6kd+2lyim0QOwcmCYwvvPKsDCqJmcegEbSHlT3lNY1FagfoQZKQn5fgjN12cm06Yli
MDRge9iAKsEZ2jp3jRhAQDClstWxJFDRaKzFXkg5NbvVxwWTGnfaTGhCtyv9ouIpVJ3RygtA5NiV
kWJxA+L2vGqE3AL23O1YEeGazYpjDSRX+aSDEddMMpJ4deKB9/KSB160GquycIJKJ9pn8UM4SMTE
jtrA4Xj1+hrRvsVgSeNPtd+PA9cUl6lRJt09xxR8tZC9xUUT/+wcJRjF/yinTB1iDXEbUPLak04q
XRBZLVHkwmB/DkzyG2Nzxoo3PWBp2U9842NUGZ1hPJ8+wWSS6BSEnlTVnHv0p4zo69RBDUrzv4D9
5p7KxIf0iMyhgEvRhBiUVreuFaM4IHcM2IJLIKGNIxtpmEPqJ+/iTtXM9qzMyliRDDsua/Kh+cDv
Udj1oILnRUF1vzQDcHdJ4VoSKBZqRZNGbyRefsaoYmeseqIVafZnuUusrSNXafdac3RgCQR0khb5
Mvnq+TSElW+glRI8o35yuw9t0jXFPoJdVbo7+vWojDrPy863+WRrn9lYllHu2h2q9zi3/tcrKRi5
aBjPkpsjbpJ3CPH8qX8NWYrcxGc0xVW9u6g/Z0x/WhhW5ei4L/cSbswkzwXvw9jtxOjj8x2yHSJP
x0xedkG+Exl/IhlVPQN6xX/n4X0ipD4EZen9xV8xjWM0TAyecbskqarNEpNnPolAA8N9HaPIrbxK
X7yR20ZY9FkiYTsboMFBpIEaJCf2T+ccDmaRhLkZSS+5YpQP/4tvjFqLKaCkeSRNx9BsdbGcLrA4
muuheR4dJvXHuULo5AIvFJjdcvz06QekFrDFkREFxnsio+yOIs8f5mSOukIcW8wIqUPUex8Gb3NY
Zu+hftWgN6aczFmj50A0KBoaf1SC2QvzBYkADRT8w5fxPeqLwiFvxogj3SzqjAUz5JDkKVnb8uqi
ATh61hIqWzOilTaUlu4CmNB7TBlFM2r96MzJ5gJwDwqfiMWctgn86snaGWtzGGsmA5ZkAYtOLY1J
EXxRuBO3Dqb9SWtY9bea0Aj9W2ZYIom6AO81yr5hVZy2pnqIpfTr8q3qviDcRtTYL4/lQl46I6u5
bVXnWp4RIqdtwoWKmLw1F8NCKjuyCZg5vgM1i6p96QnSX8wRMqL6tv77rm0I+t6bieBZbGZavYJX
1JEaVKlbwsYf4z+GMfjyZoeBfVdTeEl5Obw+uoWRICpDdmNPWC/wz2QspS82Cer78S+RxLlkl0bY
XYlEN5SLWokDPTEdwPJwJFc5wBAD+8c4l+aqnvw37PHDW8iENWJA4sdRq6IZbhmt+0K0G4qDC/8S
I2Z0a3yPW5UcimTs8tm/Re/GHx0TN31D3wwGkJCeezTUI/c/vUNGQ4RAfJ3j+JPouOtubCQfuC95
6+5o/LiQv26Mjpv/hIeD6T6Y9fr7Lk82V58yYxgNAIWsaItW8QR+s7d0aNBLKqS9Fdm/X/WZG0hv
1bwSbiEyf3UtfZdtugpB6zlMtvwu4W4R1GTerOSfN8UawDdyp8CC8C1CcfP4FxejMOVpsUSoRiAI
cxYUBrUDmWRawOGptZcMeVhaWjSlACPlKNFwvGgzlpgoGS9yrp1sQ0y/ASRoe0oYb5M9uLXlaw6m
Wv5kV04t4gTV6MLaekZ4qlp6G8z58G/BL/t4H6IVetAdAPYoWYy5ZE0T3YDUC4gnYzN5RcUoEduf
jlfVRV5VTEuRqfT8ILfvdd2Nqrm2aTsaWds45AhyC6PAtgRL7P/+PxSjlSeddRNQ5UchoC+TsDNZ
f94cRtwSo4vKQ01IpLnYJvxYkDM3GoqIjbTExsnEhNRB91M/PCmL8N3GFjOk5NsAzPQU3bespvWc
2/mu32+92VX/g+7tRfV7P019ixup0CXc3r7d66aR0C26iqo9uCR+eKsMJJ+TldwVIaYN6oWKmeg+
xdspJ/5UwZl5rAfffDUUsW4kHUmkwF0JfKyAJI8lwiBMQeHkmUj7VBPG5xHxtM2Se81GeSyPZRE6
nBEgZkKjLZ6CW1hk+an92oeqiKrYKEKV4hnXszcx9N3PZw9WIJE5+NWsu0KruvTQrgFqWtd26SM0
HHEIQPwvnh5CekPZ7QiKVBwagsH73es8KG0JC+UJKEGeb+U1ZWN9a5QE3Q4HwrmGCyD3eJudbfrm
YmqL6jAvMIs2hD2FPrRF0czeGM1hEzOV57eT9h0yN3fDNLFFCv4fnvgrriIrv7kpbLpulg72+Sie
o1d7a/e55piz7Um0Sb2k3AwMTO1KPvXBK7aiRW70waxng9sD4B4nyjA/J8F3cwJSny1cL5DhDQSy
L2aly9OKZPeWWOv9Zp71Nwh3uV7QX80gx4fMlD9ZDvvJiqyAP1uOKRLvUia7W79+MCl4GQAIUZVs
dr4JDNwA09A5RGl7JMUoD2xVlzQv0kU4hPKzs09NdLUAVxXHVSXXgoCMItCTVcHoAMrlM7b1SH4W
aJaZ2SV0n6WCIm8Hq9N+c2Cka2CzwXfNWvCPJgWE0YXEvoJxnu9dtle1OVESVNtO/rLgBq1ht3Jj
EHVDI9s3qs4EMPolBw5f/vbM/FCYv52he58sez55nk6Io1CW3qzWLlxFX9yh80pYjD0RYVOD3p2e
BVwDDGMKZgSrtP0PmER6Gqvj9WjXbqcFffNKM4yaP5K7bduOBbJg1j4wQc4RnqMPmturoyzmAP1J
Pp7ZvwsT4tFlA36MX8Bc7KzxVpmweW5vEph9Tv5GihFCOmamscxtY8k1GhgpdgK50jS7zDalgRiA
Ze8K/VrEsWB3sTE+Rg4kWlDkOx6mecU1wJkage+JSBdLYBzIK6/1BqUnKFV+b0ESdWKMl2/iSjuy
IsqgSJxHuH5aawzmtdHw69Wdx1qPDfemH2KPrVnCs3/BCsrqm6gH1jQ6UyHp4NoMaKdXlK259xlR
QNy99/LM9kJultWV5yCO9d8dEi8VljEIVPLnJ4sIwPpi+HyA/yy1f3zaCedjdwoF0kFYrXm7mPhY
fGhC320Lgvxc5Iv013bzsseWPsH2ugBrD1n54HcqPG565ZDFkcuSqSPDUMIj6y8F2Kq/3dkUIkDb
y3RCuu2RHSX8q3DmwQoQ+uRG393hZezOCxVAm323r0BdZc0sSPXM9/vg5/gRg+DCCHBVuQfEsvZt
2DXP2VL0BOhjOBm8Fm639eUzvB+yyH/7rXTtGx+NI6K5AcGGsqUyr6puTrkwFfPx6AGVVyv95/4i
oA1ML35kZxwYuho1kGNH7djwSFKviDwy9HVtCgPAEQhP+HwtjzFWPuVHXE4rXVLHi7+AsdCrLNkf
RFeTi7fTHTD8e53hBw5sgwtriZmaG+LAh4wM6rise+MH+fNEsuku2qsGoF+taSaA/2s0HjSKlDfb
i3GwiC05bUqQdFuC/n/zyHJY8AwbzvULaQTzak+kgkvIeiSZhywHHUW0N7EnkkF7OPd3FZbCHmY+
WQbrbDx7fFcii6/YV26DhsPtF9zSLKHUNJxKDupNF/tNOS0ljFnklqQqY5KQrvWABUj5IE6jyzlW
UZZGuYI61RGGYYyPrpyxJ3x/1lNaYs7nKsjV1n4cZaSgd9Rh0QnEoWD7B+jcYwlTheVcQBR63+xk
XzCi2kpo6Vdm0SlNG80BMAM8eLlnTFuRUWD5r1EnjvnMDjCxbTq02rD3hPj+qNoa3Gs7V4pgpjE8
2kzsuxWGUzo5aYGeuFK3tGfF+79JyZhpiDLihYIy8SpaOGERkFbA648xQV3Mk81ymLSQJI+8W+4I
zAHqUiM2BgVMOgjx6xTVoRQr0VrgE/+Q2/mBIfqkJd3bsiKGWSBQ/aEt/APArd5qI45H7oaWMjvS
stGSe5TvG4S78ZlUt+yRREoI9xFlAHD7MPeMYOo7HER4uAj81A1U6Yoord/19dZrbZSHKtEsVjRL
6syQROWkdf5L4uYdOCpPwSMPqQntZa/Wftt9me4J0jonXlokKWzCCbhJBw5DEFXJRvJ6KbEMBoU7
sNpB/H09b9KTeotAszjwl86lIBZhfyJ3c6GOKAEsud/nvZOjn/n7bJTKgiFdZVC5hd4eZIVAlGsk
22G8j8GJY+yUvf9+C4B5SA9Ruw7HoXybhioNefnRsws6RNpUD7gqbpwdTXwyfpzPny4bix/Ae8vd
p9GZXkdWW82hueSHIUZtCwEj1IKtqysSkRb0W1SSol9x04ngVgbU/TVeuhHfPEONtSiLtuuG3r5x
jvUjCNZ12rSago7tYAdEGCEFkdyio+CFIRX0dhH1jjG3jZON9FkfW2sml3JNJJhnn6SNhjjGZlSO
wg/7FVjt1r4KbdTPQEFYs/vTdMd1Pyo42ENGoQedLCi/KNdOr2Amhz/npr/RqP+WXas8WPjEh+yo
CpXnE7XAyH6+Tktnmv58HRv/XMLm50D3ezK6Jlt4uFBJNAt/mkHo0xTkoyTHzMLXtf/eD+NJKIIz
3MNyMMfOGHqEhI/b9prLRPrBOYe8i+sajUr0P2Hesmu1W4ymLyORs5dAGMkwILrJ4D1Wg911o/zd
dQVeRe7Tq72kOvdfBz/33Fmgy4f33vLhoAhjSZwsPf7kY5Ipj5CIxCflALIeslxFiLPsQHl3EWW9
wXKe/Wraxy8uQDr97iecaatkH5l+hXBujNS7mV4zLNCwEhOLYSbAZR32aAYhTZzMslEtsbM/7Ise
vIvDQAoIrzZB0UxXfETyNAobUXUhKVmRTzKGdAmfWUh8QKqBvflfr/N9HgNdPmumMhtr0F6VuAuu
C8wgZ9Vkhh8ADVZN/SB3L7U5C+fc9wdcc4P74tV/XjcuQyK7a2uWZvNGlZHU6qlrzgEvfVP3+gU3
tIM20KAc/1n2+zcqyQm8gbtsnqjQClzNOS5SXZyMk3/CZVjljje9RrpaOkn2DvpHLK348em1LWGW
+B/t5E7nGQlgvHHrAxkZayoFA1nmq62RVkVedtmo2iDyr0+aTO4rL2TKTt2v2kKHkaRM1cvh2yJQ
zOUOkrErcWJ8DXXR6xd/3LuGKh5x3e/7/imyq6qH9mQIqMLuHRZh9DTbx3TJMBgqtMddcM3ptiRC
05HHV9KhEcPzMeRO6r9oBH+XyEfvNJdpaqhga4Vtvf8HAcZVGmk2fDoqfUCm7I3Wow8Gl0/IpHVi
+YyFgfpeaoIbsqRnyQbsoE38ZdilDbqNH1f2U/X9kmeVH2NDOpqb5gYDz4jyhMX8NBHzDNOvn/y3
BXHPhZW6njdwpacRx0O6e4ZfYCf4c5JTx0qTwKh2CwZPSDSYVQ1v5uqeAuE94aJt+Ym9r3NQ19/x
EY7lVtdIazTh4TPAvusn0zRmEWC/W+3u1W7Fb2vMYIi6xhzFJVW2N5ymdJWVXaZIw6bDISkTYY19
ke6DRkyQK+LVKK20pqfyUpTgpIXjNi06B6LFOurRNxibqyk7YsXUp3V8lXId7H0PZJcT4nmf9mNi
5027iDViIff9lboo8ywGORiHPb07cQWMQZT1eY63VxzW378VzSJep4TLzzoi4edvDWIYfBTU6be5
YHuOCdKdSYucjfNRjepb1LYnaDe/A4A8rFZbvHvubn0NCKHQ7Gbk1z0bYKmKIosi+ZtY1F4Zakki
NZy7uO+Iv1zIyJq5rmDuSZvp9I1X8/pX2OQnl/SkH4NMIM5OYk2L4GzVawfZ3Q3/TLLBl7ec3Ttc
87pcWyxWUPCk0cgmf67YuRwh1Z77L/uw3KzPIXNrJxWriyjVAx/tHlkw58tMWaKMNY4bDKEXy1Ta
BYvrp0IuDZnVXa0snwilV1BVtg1ePhbTq5ivcY3UdxUGGtB3Op78+zAFZW4EZTHQJFlZE4EkybYK
LcXNW86ld9UCJo1F6d79znxlvrtZmWhfDOSGppwzbakC6E0IaG0l7dwm9M/HiBJ3oLIHCp8rJ31s
Stt1DMTpZdXIA1p+wlpWjxE0QvcbtucmneGQexbDtgqAaKcKByGvjcNvAYPORiqcrrpxjAckDvud
ck5ep3bx2YrHeKFMNTPX1swGoaDpHhhJjglA4CmDLWq7Gnie3wwjOZeziuAz5TE+VL7uz4HlJdcS
m6U9VZqjzSmKIefFQLRBrukAr8rg/CgNtbPDAUBLqZXzrnuj4+4g50xylHlXePw9NOX5gSqGPjQZ
C/Hu3VRwX1wCHEp5bzIxB0hsNETVNIDNsUzJSh/AAY/ARfQQRVEASv/smxGUvGoQhz19Q26x4amo
a6WJyvmGCcS3FH64UP/zJljYqI/7l3Qc+MHyTsJyExComjzSkUfxj9LphPcg09jbiGgVUrJ8SG31
7VA5WFgtGfRu2GxnldiKRO1fyzwgLiLcJHzCi0Qvtxs92ssaC+LbuaQRsmEzsjNHQLOQpHjKm/pp
Qe8xV0TKvcTr0lI5k1KywVMwSIUxy6RztofKHqoitg5kSAHJeFvDkTUbCIGV0opta65bmPPRT48H
SC0ynMPoZ3+DUJS9AawiT8IGr9KuCtO1g8AYR0YNB9a3palmRESgehE9Nfm+71JzC5S9RDmGU8dr
Iz83FBkeqo33TBmc4+oJzi029LRqy0vPlTYdLrUdqnDD/rGWZELYBT1Gm4F3QYvrQRccHFjX2RVC
2C1UDrOv8trSsMRqNEHNotr2JxxLUjFqshWYQ8fQaZhxoa4aB301SNnhigpKL4RnLwG6UL80mrWU
CD/fpG2RNcEW3JaRGs8h9Y4Sh3gucIwRW2VZzZbSRQpP/KcTkCNiutmV3Zu9WSjtXiOWyCoZDxVY
HSBuwu+fTnKkO6go3cuFv/O07YBSb2VnTr3+XTluEeM/A4KYY7lF7nFYrqCAmce5F+gg3n6rpmtO
zQnKNYkARaFcPqthIR9oD9ge+qHTkir1ZohUeBjdoPOyws48apyStr2n/aSfZi//rETQPXklDE46
0Y4LqUhj2dVSZ9CH8MQ94CKcx0smOg3YXPRnK8mkREzhsgQ5JMcE91qts+7Q+2N8QQ0gArHZxDrt
xPn3RmAHC1oRKHYWD9V0iWPvMCYgghhF68cMV3v3ldACecBZAX0ap/foPsgjJZsnqvIQaosIuak0
8MVE2DKk1td/sebnXn2PkIQEvMnKe6t2mP6dDJHijkPQ/CLfXscex/aB8xc40fgeLumny9XKALCa
YET52QHPzbsUqtyoXjomSv+gJrdvRkluiCgJ7oMwZ/0LR/44g2WfsoAITXIoCVrMAvIcLSz7hven
MuIkAZM3VXdamBJRipdqMFnKCPsKsAZ7mPCMv1TIO92Cd0MIWnG5R2VvSNlf4yiGqV6Fnhu86kUp
+6Pa47WYL1pRBRj9SOldD2ffjd50tUKuYOEeA9x1YuTwnO+uSkRdf9Nzq7ImtmN7u9vCeAUCahGC
xMaIr5M6AmqoW4MkjjI3wID5Mpd6jRg3Sw6sSBlGHPGPm2x3WWR2L7+IJQuvfaLhPoH42HaakLAj
haOPNnnPQKWloa2UlKqb4Gqc7OxmpWlUFkwAc748A4Nqsp3zcv87F0I2bd01dVcIJ5MxWcdkGAIQ
iHY7hb8DlSPP2Eq2Du7s3IsR1oRucOxZGKwycnMU+qLhkoLvEGPA4j3yraICmL8dddlPvH7Byo38
jF1ud5suwI4bgSHveva0FxEcxvg3yeMjxJUAWeqqIqm3L/CSt57EMyAz0RX95INlfoGkAIl/xQCg
faTutvjYm64zVPDkv2BUk+VmqP+I/Wx4sgGJT10opUlVki97PT8Ngx/dCShwRRu/1+S08CejPQRy
QtBqcxboN229xE/8ZyLixHs9LP0Q9OFPQxkPeRDsJd1TfXwkqnPj38SfTFrvxSmlf1Cr4IRbk5Jk
T/VsSTuotNoRzaKmnFr9g+kfv0pGKqgvHrvMi6qRmRUdw75DenS/fE3DDt+Y3yNg1Hg1ank6Bs8+
AG/DPNdifo0Wr4brxNgeQK4fjfA81MoWeno6OWZfE82PqcbOFjxukkUz4wVCu87Lu0COokmUUlac
+FcPRSeeXn1GYpQEdgWnLcELFW5JBymVlDx11gm5dLCQrndx7f4iIH0oOsjEP3OnpCqLNumOMtWA
S9GlYw6V95XErJLVmc7kyPVLEx4P/F2GhF0rB/8XC9orx9O8m57gPHpVLiOZ68NcDqbW9C4qg6fT
Gb8bCPW8y3XYan+zmVIkNQ4qerXc4LxZdCaC1BaGkxsKsv1Lhs4WTBJB/akTorTtzvSdfJI3bXyl
tJYYejTMlKPMRIePi1fLW3jr4roVNFD8mU5Ah88K6qlAd5p95wQDkkr9/rLnxlT9ullmB71RsLkd
sneC3ltL2soB7caqszzdcBMq8PJpc9wZK6LApwR3OTM4DHpktLsoMfWtrrXNfx/l1zImrSrdMB9N
IPaGJtupEAK+yVdtk59wo/NAkHgEzsEGppC6p7Zx8srmJkuKYgDEHEWSqCYXm2JtjdraLi1JsHwL
BClEWb6gQNhwgI7O3FJr4fnlnqpZot4eFRushh54aUxvaINa3qHe3/wt2gecLBagY819Fyk2Xox2
ROgTIQKYgQHx1XxNaqFiUzY1AD9K9+5Hivzk2NgL8/PBaLdL0F/3yHiLr8ejbx2OBHAd7x7/lEq5
Hl45YYJNs+jsG05se6Lz/63FyAeD+IV9tWrnA109UDzY2O2sEIVUsnQoiLUKKrLUiGxnsLD7ty+W
3Cum5kN0xqRSgyp7eZpQB9Dxi3e2B/qfk1ROH9LVPZK5eA7B3wbRD6uw3/SOgQ201iedE18Wc4uU
KRJ//YuYTU0GyBbTBLQUJWJUEubP8EVQ72BUPWFtWwx3uBXw9HW5blIlAi5M6g/LjPfag6r8fhlG
GUPKDgJ+2vHrgGhEMztMIcNF2hyq2SZegr6+pAXwGusRAwvcX+WvSH8JY5z1tVaH3L5jBL+WBwOq
gB6XTUpSzK3wpkTvKTEAKwQBHU62A+gsqqjh7dNETqQCKTxj6D/SfL1qJ8qZXPFyY+JpTCBdkoRK
6B3VP3X+t6zqZU2b7M3IBPU2GUEThf0N57w7Ehpk1IUDAKn7ALndhcPkpmSQaoMi9XorCh3hPIcV
xi62fFd3zfKCvqvo6vOQTfTSwiWXDx094XGLfs8wL8/HiZbvcpy2DYKk6XRhN1dLNTG8KeYwiwDt
14NjqnnovyyuaPWQoxI4hdFvmLmr2x9Jo1LALVgKsKYCjzMb1T4+vJ10RrKTM6bYvyU0nVJVjVIF
NOydUfFqMBNzSOoS+rMCci5hjwCMtb47Bj3+S53d+TAptULnhF80gpKq1ZqqQ+nNGDejTRfUzTqd
SToIdY0WS9C0WXoEDwSBep09PDfbS+CvrlEdvM2cmDT9EHnynUP92YdbSQeU719p0UW9wcDNw/9k
NXgZc+idPZkRBc4bOn+29d+bRGY9C1NHHkCkEm6vDzIA/W2mafdgyE9/XuAk5DNYKkUvpeip2uqK
ISWkoyTnpQ+0JQz2+9iUhNBRSiawhv2mD6rhdAfmj0Qoz1Rc7cGk1LsSi4s1TUjjxluJFp8zJxfz
Ukg1/wNBR72ZFIbOY9nCSdPebbdgRP/jHgkA9P2TKuBOD3kRExK+Z8TBoHbLpowvvu9IJYGbEUFg
Pm9VFlBzFJx0QpD/rqmG6YeoOFZIG3TACdtapAyn4QmDq/9x+aZS0m9tUuuDOSanjf5Cs5AUzRfZ
oERAHBaQFsLti8VpRK/Sk/FPDHW6mGR02dq6rb8DvbcrlxodTXgSHmx3ZkU8U4nz65fV+mgmGEml
N6dnIPZhV5PDHZINSZAL6M35YXo2s4y6arpQeJVupS/ODBKAG+Sc5Ckj8QuBV0FgHBRFBlPf+oZm
/lZw5oCgRUTNtVC0IehPVn2Vxn3xkP06J/DQuktuSP2lEVCJCmyounP+IC3GlCYYZuiL6g5owg+C
6pMnMoHGZuJnL1iV0P6W3mqm4IJHfvmt6XoFl9FowVyzmOoVxMdZ/kqre9ar0kUNr3fHBp5BhPKb
09721Aebl5cJva3dMhuFuEOeGWKp+MkWJc+t7NPZJLaDNmhz7eWTgecq9YDl6lF+fs45XQRImKCY
AOabQOnqPoFReTuhR3hkI+GLucmkD3LpH2DMFo/J8Hwf0UAn9O6RbH0Tpp/Uw6BZJ/OO0CEk5PHI
MdrswJmKvgtPOcN8hFz2QK9wCKnkUvRKTzoX1l5L8NQnAZ/BQ5UxOS7ahzHodfJEMsvHN0/8JCNn
3g1v81DU9pp6SzZT2PqmmUG9sFp1xU6ro4SY+s6bc9EZfIHaX6mm7jD6EmdrY447ZX7MNEdzapK+
NbiBUiKM4nkJFy1QUlSg5umPAFpsDTVyPP1J2vnoMGJHZAyLoEHIHC3UDHqjNS8SgKkUThy+bvXq
Oa8N9dhexOLBMsMeVpbNxYr64mHUwE8fHfuT1f9KkEai6Wiq7aA5zBBdfXAFXcbBHK7ai/iK5oyw
A4HXrWXQTAAWO8zMb6JZSsvqnpAGOztAf4WbTGSsO9ymjSC+/Lv+6hns0TJKh1LiepUX7Crnexg3
Q/e/wy+IL3KvMkF0oMa0IXf+UYBplGHCNIv6pMFa3aqz2kiNFv7OFA/76Mtl1m6ustxasqkgpHQT
ktXqCGDVCYEaHzu4R+Nk+mQC/S7jIK/1ZwnF5tt+54EklAB/c+OQSNjdGNXmRRIkpjeMJLM50OMn
L3QcXIjO+zQ2aT4nGTBJPVKJxAWA1vEdmB6+QEXj+l33Yw2qE8/x9MDJ3GlUHpIw5jdgXlgKS3SI
uKU0CGnFvqSruFRuCTx+CF7oaArxyyqzw5NEgXhbAE+0viQ58eQHppQ3Z8yG2umHepcDNvGRM3oU
/LBkOrvnFWlF/nHRnUswVJDlHPALESK9TI2RNcO9FQShnx+jbIUeTod5F1/YHm8XDytGD1ZffMBY
fCfy4ngk+YZpvl2bqq4cOLlsw6EgQpEOLwCMF6IW137uxxdErxN86WnJs/2+bKQ6ylaJDvNvhWtg
IStdUKr+xJK0ThZCzmSFNZXXUjRJFu8zfXAZ4wekwV/FKU4T5l3q+EvYBkRbjWIcXxb8tmW82fgH
M/XuJQH+5aiQYIWlebNOH91ORK+qWt2PcgCmxOy6ezM/ZJlqDT8XoMnordVpf0r/0LvYZP4CCMtF
YWtQCf1/D5V0E2CAFjRf71rnK+L/qk0jmvyIX0MQZHSFL98GE1ErPSUxbnOEl3JzZonbPSZNGplB
0l6V/BowhSCrBFho7FB8bizmrrdsdlkx0SkM/9ctM5xi+ecktAbdL+Kl51tNorfIvXNzm20xAdOC
e9ADcfRtAzqDOkieDCNrYRka/vQD/T7TQcYh9KHKixT/oPfYLRWm8BMHN1iwqivut+uXOP4TLegX
BwwfjD6jFgeyq8l84S+lo+1sgzrRnvUfMp1BlDrRjXnmIlthRkxEvQVnXG4THsrXRblTcMiBX/mR
XrXiJOvuz4jN61G/XxZyeSOblfP3BE/GCRYhdntwhtRXCTh5FJEWkG9xmnqq90CXyWIMs7esfCzZ
H46HhTBb+Wc14fRDTZHaFS40iFGMG5EZEh6wV+6amY9S+5DshbctS8kvUwqm/V9cLhWihwltHgGd
9b5oktajAqZm9wdjjU40NZM5arFSOMBYV4/HqimjVRvR4EGFM67nYWXxYiNPJl+vDfbVZf3NLe6k
dGqzpVZXIRFY5nAACQQjezicrXszSbnx1rv+6eMFj+kQjuyraQMWZG2LdSb619qJB7q2T64Z+iu3
Lw34xHrmA+/KuLffPv6aGBGFZN5bBUboyr/xrrSs7OnDon9VysXEhNzPH6aWGebRB1hPNHZAIz1u
YxlVpD5lxoH3dB0xmXwjJUtX1Sbjcp/BOb+6SMClXm/EnIi0N4EtVNbi9xBfDzqH6ZTEak2UD3pQ
M/y25okSQ4+bvlZ3zXUveZhXbmKTDj3MuZcnF0yeTusrv1NSxvWxa8m1yFejhqbZfN0925SOOmH3
iVFz8/0iAvecLF2YNeMbSKU8uLmVnJpFDlsljigLugBrHKcjaxY4I6MT3DJoXUPORSEtcsAAngdl
25uRjwrIEDCow95avWb8vLwOuiXGwC/Q9fmvIgygtPR/FTdBgSdsaPBJoTj4tCMUcvQ9QcMug/Q+
7uh5Hv2uQYPznXBGAsrcQuvUT0oLWp2li/Kgghb5AlUykGWdiKZ4/oQfzpXY7Xmt/c/z5BXwOvHm
LlwWnpax65Z3KdtvYckpm/+5r4pGVzqDLJH6p7ay/mtefH9mxi2jfSh0tqNvZrkRwv9KOrXH/uK0
kpwm2VHF1yT4dK5OPC9lyghk7vtILl0vohOezozTPE1M6+ka8tf3Epi+MaovykNGWO0O6haa/SAV
IKrwriyXJUMFDCcIuRb1S7JQcL9bvm6P+KE+TfPIx4o5RHCd0YqSI3UL2DJFZYGtDX6MIWUm7kQ6
f/oCR7v7/hh7EjJK6WDkjmWrKEVgn5EglYUTk+O5Zq/M8I+ZWwfSLII3vCt9J91gGogvMMZI8JI7
wauJYbFCMn5RIml2PPZ0oCFJGd58oWCODiDd7IyxoZuWeVc1uMQUiQgIfzjXvjI2ILgfLu5FvSt3
Z5phPy6xzJwjaG3deQI8NU/XjwXJ3Dc/3ixvCKYrZIxvNf7brGUC6UuIJbgabrftqLddDT46jToZ
/i67EX6qXXI7zdCs52XIk3xyK4WZQ7t950eS72EcNgGQGDWag1kEpOWnnGpJvNayiO6yupIb54WU
fifluvsC30bjDAy6txyjFmab45SPy97qskIH82fBWIwKWnExgR/rq2cTaDi/4lD85T1V5gUwFt+z
3LanwjY8C2etJ/H4qae/4UCdMYJtGLROavwZk6Hrwu4ccdaN984JABUjBVhNsEvg9OzjhvCB6pf+
Pqtsa2Z+pyu8QCckSpuoYL9li2NHiCqqod4IG8s23FeDYMgSoOLnoHE+PPwnIn98TgOxiKNG9nCi
kCU0Nf1FzpMMk2I2YwAhTVyWRU95EQ37bVoleSrXterJKBwwDqfkRcoMuzwUAvSoLaCwJSBLGcI5
3m0tC5/aVamPb0imtI/vLQcXQMenTWhHWAWX26STKTEEiBFZzLYtyq6oMa6j95R+bZZwn/ZprCVw
r0NHQj/x3K/Gq56Mg4ecGPgXqcAm9Z6FRBd8CFhjXKO2FuGPuCF43OV4fShY0U2DR8PYQT0mo+sF
t716bBbMOym+4VMj12usZx4PCYqJWEa9mEGU2RbiwkbJZ/KSLW3Y/JjqEHuG2vstBl1ypiS9D47F
pfbZ9a6Vnh9lWpvZ4qxm5DHfMfWLZRl16JfxT1IShXKG6bdfHOBazcZxtLT02CAxKtxs/YgFVYLb
uzmevDJcCZP5vl8YvXbaZPhWpSEzEW/RZ2kMbtSXaseVRwtTUGWWpptH9L58bApeCpds5z5B80OE
6fp1ZRuR2IAzDSL5lKrXVxbse3moHrf/GNe5aUDmKpucv9xt7jdPGtTTnocHFutq0muKJ3Lq/EM/
av04+Q3Ttf3uHmW6+2Dt24/hvHYwFQvQ8EB1v4B+zkyZUbkRlVk4bGAg8DOuw1oBS/McqJaU3D/q
AVr8hUo3EX2vpf3DQxFoHsa8Nr6qKQK4AzYYe+oK0dNs1484XDJObdwmyYzYE95GTeDS5lCd+4s1
z0exm0p82kfdbxzwOg8SvO3LN8RjM32E9V6X8+fy9MlVJ0otAAv4VnKYKwE+IrX4ZwBFPamg7tME
sewyJS98XCVDXN1H0/dVH71ewwTKDTaNU92NSlRNfDxrwuoRyfYwpG/LC/6Qdlppwhd+Pe0xNy7j
tpSn5XhPZVfDHTGyUc19C7jmhOdKWg/BQQFINgencoOOTvW4jmOoueOGtmDhjJkBTswW9R/iXFox
IzhRCvcGmIAUyMpw+sL2a+sY+IkUi2Kq2r6j33G+j4D+Qya0ucXZFldMPh4lBLba9kGyGU+zQIEI
kbQ9YCA3WOI1LcQuTj8WPE+hO1r7OgIunoANbsJqnNV5JtWJ2u2OJ+466tRU/cUtbI1vHCaBUiBB
EjLMmhNeot9p9+xzL3l/nW1x3PQ1Dy5eaw/L9MWe4z4bKZxHCiKgadsksj7RS9zzhi99u+EN4Omc
R4NPweSX8VhOkS4j1j0rImmEjaSXOt2q/OQ5uHSIhZxf0hfJqeNRw21nvY+RK22AzIpNPPFNfOoO
zKnDUbyjzUHEIkXz1UPPWmEeA3GjDwyesp/s22C497/rOFm5notUHGNJLdA0Rhvn7DnA++v0rUN9
s1XRm1kew3kOgj1Qn21tw4fCOXkhP7B30qf9UK51bFBVlb8ziNKpB9fxodyxr7wCwS9Xg4WpLpZL
gKw2F2t8wVSeVJFGj5UqKVJVZ7OTC+LLqDJ5MhrSGS1p2B16k+KKoJmk9FUFIKWwGJ2laED+hk5w
m+u/TJQwVZVchfVoCz0qkKl26NcqLclTK6FdzRw4aGJd8V7ktp9+TyPgiKIkwspuqoK0CE8jXTH9
NfHmK19STrdGFgT/Y6XsLoo72eKzrQRFsqu5DGi3RZ/CGEz7q//E0celJqh7WOiLmwyyLqEOApDG
zpLKFY7Nw0BBG15HX9AATonKZElb4IE9pqOEnJf68juA7VnjCJeSdH3i2HdiyFFdr68tFY2HzhmR
Tvxv7MEAyGhLxfnWFAFsZjCL19tMtEp7c5qV0MW7Pw7sEWACm5zoQU8Wc3bDgiQxiTNZcWm3PF90
LEPUNcq1lJPY/fmKHFK0NHpBwhuVZrdadoOq0oUAY/BTvXacAieeqixXZ9tDGUyOkh77pIHLamRS
QUgGvaKRucY7L/rvSQuTm9FJs35eyNvFVs9ulBQURPxwEz9cPDnerO5Z38hcgT3xwOzQLa8huuZL
MoVrrZkLb3mT9ar2LdcTpD9ODw+GyhFcNcFdthPgE2zZLmDLkWN60ozCLuEtrgfHUvcqHoQmGV7L
NAlKKxqFcBIZcK1RqrekD/pd1DsO52cGSrG1JZV0KsG88praSJAdXVeJJFxqLjLLpzJPs7lPNyau
fSqei9FKjZCgU75J6RDebzioOFQrt7XAXZyNQmK+b6CtgED917QQJLYvuj98qv5bNb2LHJKd2IPE
4elCm+bQni+ggq2GHs7QYrh1eVFigUSZGJtmngsM6NhO+JVTPecm4Sc1BI7WuOaLPHQ2tZXIoKom
6a5QRA4sKf6fHd/6T+O0q+4RFl2VJhgCCrcWDVLsKVYhcP9NQWwZwRrgoCLIXHmx2vKBB3tXe4XF
TMrDXG3d17Sx43ouO9eO4uaM1RheDztyyTp0uoYmS1JFs22g/DWWHotWSy2TI656eSltf2JRHktY
Sa5YpPsSeE7+omLQdr+t5LVxhBAMIQnDgpG/GKEhFJbYlJlGBq0h50Qn3aIFYO45PyWw2xpUC7/v
TZzu4vpKoBwErYnJkR9aZI2tUosyo2VG3blOikPfUV11TwnZQ8OLi6W3Qr/g8i4n0ueO4rEfDAOL
iIlircIQk+ZRITPgtGgZOGLqpil1ss+ISm4h6SsgDgbhorAs6OuGwl4m1IXjJI7S9sm1Ej2U/nCm
7idAAPBSPiw6OXCuqlG8DqhBwhYm+IUKOISucCQuYM9ncMEtCOOmh7Ww6fzfGxrKmGo3B0wwshSE
tH23evLKJnXOhfMwwFMsnWMMUUpTj991LZaWl7o4eSRAjoVxGl13wUjSiQOTUtO22MMJroe8Xc2Z
yItu13vnnhTcsOUa1OMbC0TxBtUZ3Ihk/7j2F97Xyq/kBHbME3afa5azkXkPNOgH9JG7C8LLwgOu
S8xeLFA3SiUJCjjVclPTdi7zHFukDmoEfoE5MzVDdE6ijUwF90KlkoZzh8Q0nL1mya+7pC6TvoTy
OnVw494yoeoUmNZ+OwspXniCeWzLu1C/8IVqtgTt5d3YzPrI+u82Rn7RUuiFdliXfoy+wPPbKVje
IOGgAvI5S0o3je2uE1Hnt2/OGdBGtTRYN2L73XzHEQx3HX7jaKfivWJtSycU6bDx6zWd+iSCwOpP
LZcyr0mC5PLS/3hsnfSBMs26TN8Zafw1TKl0nhwdZAyWjhofoKqtNrNXxszIhGgCH0QiIwbjNcVX
ExxcRKsfRyHkwgAk7QalyaTl75lIB2vO+IV6JBKh+8cz0Olzlx/Flc7dSoZo8Gah1i9aeAoE+wS3
eCqnpGLT2DADxGM81jKkKBR+Lqvh0Yht1rHBger9w2Ke2/2abKPuOL90fCDoa/Di/cYV4ld6JCpS
aPAIhbFzWzGT90kqip1X4cy4Xau2/CzQXRFtaxHXt4Iz7eGy35OG3NpKmMkBfKoNpO8tVIhkhZS+
a6YmVtEbHUCNIKCCDuUf3dNcnCQ0zkeZguwR6OT/I+33lYV7HwmqkzNhh5kRNOgsNSHiQX1bS18g
TFF6l9DAobsD9QBOq/FDzclLzfJd3MwpLsDInE0viLU5O6+ydrBb/KgPpJ78xxbYFv2z+P0OeX9j
4FuwxtWPtMnr4A741o4eMxBX+kx1j3pgxBEe1tOrVTBtdJS/iDE0Gv1hU0TnJMRoPqcsZif4M97o
7SZ5a6FRjx9mGP53yzLC8JbAc46h5jjRvZiyqnlCpED9cP6cUGIXwmRkLspog1jXRvSCEr99tCa8
JzQtgOZu/uA9n+KtWTTtouMqBXZt3NsuDHgzzFefBAss22LZdy+YDaRRK8HI2oVWoKhQt/GNE0yu
sJ//u0BzLLCrnfJLnJ2Y2ZMh+MDqYYPMALcGyXvueZi6F6osRPrfL1BmScXpajxq0v4Yrxk6pM9w
wo1XG25wjs3bNOUufbWfIrY+Ce+dcpUVcWbDLIWznyglKbYfhekjJe/KsSP5J8zEhpwYOs5HQ48e
kUgXo3m/rgABbcwjX/DikKKKCSR/1JDQdVybydV/lBgnDNsx+ZWSWCjKYBGG8ouGeLvg+S7//xW3
A9Z5i0QBcN/YnFPqLjLYrSZbyBgp9OvxPDWaBg6RXqW2S8zafo41FzaxWghBIPrjHRju9KYXJ2ah
gcRqjOWER7s+sDOdGYAx2IDuUpCyu82nzdOAlT2vx5o9YqZLyDZu4FMaKOFLcOmVroV6MKm4zGQM
0VCPHffYJAFtFZzRhCLxKUa43ZYfnH5XghS3Yoyq7N+90TrwvKvhQJLHFUs2gRRBF0Qrgb+sVK1R
17VXnir66SjEdoWwhswrdU7OW6DHKQVrMbzotFhXNgUGKezH8k0jL/c60uQhT4na7iBFEHdDFyIo
C8vGkjF16Xb4eZLxvQ6UqJo32i1zlffsq3Z4bHuCbbcMA1z4em7uiUyrH0D/MJtuWFptRyzDtV6x
lCzK7lsNtrvLzcQ4n7WWM5WDWEtrhYPACNT3bMx91ciaH4kG96Xu8hgwvozWJZDVb3H2JvHqd5ND
fDbTm/cnqc2CU6tX4nE0z7xS87tAzA2yISM3FmfXmTjU+VDNouWAmGxdpkJYjP5XpU95z5jr6KDu
iCgjRK1sQEe1OxZ4jTyjLiE/cJvk9XM6mjlG3RCb9CLQ5drX67GClXKZAcsyRwP04jasogPI7+dr
SKguYucmsDnyBGdnEqNVCnLdq2zrV7Ftu5uqd46t4b4gR9sl53/qN9FyrILPg+VCicNeK+gEuJWn
2OgiKOm+vfnwusInxDTEMcX5Qa1MQ4d6FrOdNC3FBbjDvAsA9IOExogblqVfxjHzz3BFfVuQjUTo
Hwhw4zDDlY7Z9B5yoSKn3seVwqy7ukw7wiG+T3uyrdlHWtDLBNmzQHSDybw122YUzCy7qU5IBUSW
uN+LrznWN4W3PCvNgFR/zxKPjK503SyOEITV20ZdsJQuZLbjw4xpmAEGlJ6n8bjC5r5Yrh1ac+OV
LY8Y6fJDCjazATJidcOWli+DUgycrFGlT714x2vKU2W7lIre3gUjEf9MV9FnGMZc+Ad0x3IF8o1V
Ur1DFYsYLs0CCf7ZADia1cHjYaQGYFawoTdIfbWbEZajRpkQZx59anCRBIGzroZ4gW5Wht2CATq/
n0G0yUiPma0GK5r6t4pfSYvg0oHWyJ/VovOJw5lzfLv6Sh5ih3/Qna4ek/DFu2OzOBqTnng3XlMH
Z5VWoyWyG/JyW8aeByhdBOi0fWPMI0rI/S+c1mHPS1vmOZvNBphUf3mDbe4IUWhFvEZfD6P/+J78
eMf+erACBMlgEZBkAx2sYzPdvHh2PSI70fU2JOzkNWZivLDx3qWmL8vRAUXGI7BS7t+yXPnaeb+V
0e3/NEJnCDKYzG/PX2TejsjeG1RGh8qqEhQMxHD4ttjC00In0Vm3Fl6TZNQPpXCQsv12/t2/b3Yl
h5RYaCC11YTUtjXKgunZmo8fbkl24KmtU5D6zo2X0vsFG+tNLcwgHo5JSTUiPTUZsH5UA7H/KQLs
o2OI0q9XnsMnaI5MZOq4tbpFxOjqcdKajbU4QhrrbtHaZDtF0nqOosRgXYzcRx4JgKiGy4uM1PqA
51UodS7M1HBPrA/6l8ST71jp1E4mTQnaEYiYVTGPXmHzawn6gUnCzQ2WAk+mTHxY2QH3r54jZChP
LB8LAWOckiWJXx3ICdC5pR8QRhj9NjLqpYigL1GWDKk0E0wgv7Jd/ig7S7v/EAjcijHvKgFj+Zzq
Vi5yM7Knh/XTHUdljRw6AQ==
`pragma protect end_protected
module DVI_TX_Top (
  I_rst_n,
  I_rgb_clk,
  I_rgb_vs,
  I_rgb_hs,
  I_rgb_de,
  I_rgb_r,
  I_rgb_g,
  I_rgb_b,
  O_tmds_clk_p,
  O_tmds_clk_n,
  O_tmds_data_p,
  O_tmds_data_n
)
;
input I_rst_n;
input I_rgb_clk;
input I_rgb_vs;
input I_rgb_hs;
input I_rgb_de;
input [7:0] I_rgb_r;
input [7:0] I_rgb_g;
input [7:0] I_rgb_b;
output O_tmds_clk_p;
output O_tmds_clk_n;
output [2:0] O_tmds_data_p;
output [2:0] O_tmds_data_n;
wire VCC;
wire GND;
  \~rgb2dvi.DVI_TX_Top  rgb2dvi_inst (
    .I_rgb_clk(I_rgb_clk),
    .I_rst_n(I_rst_n),
    .I_rgb_de(I_rgb_de),
    .I_rgb_vs(I_rgb_vs),
    .I_rgb_hs(I_rgb_hs),
    .I_rgb_r(I_rgb_r[7:0]),
    .I_rgb_g(I_rgb_g[7:0]),
    .I_rgb_b(I_rgb_b[7:0]),
    .O_tmds_clk_p(O_tmds_clk_p),
    .O_tmds_clk_n(O_tmds_clk_n),
    .O_tmds_data_p(O_tmds_data_p[2:0]),
    .O_tmds_data_n(O_tmds_data_n[2:0])
);
  VCC VCC_cZ (
    .V(VCC)
);
  GND GND_cZ (
    .G(GND)
);
  GSR GSR (
    .GSRI(VCC) 
);
endmodule /* DVI_TX_Top */
//
//Written by GowinSynthesis
//Product Version "GowinSynthesis V1.9.7.02Beta"
//Thu Feb 25 16:22:41 2021

//Source file index table:
//file0 "\D:/Gowin/Gowin_V1.9.7.02Beta/IDE/ipcore/DVI_TX/data/dvi_tx_top.v"
//file1 "\D:/Gowin/Gowin_V1.9.7.02Beta/IDE/ipcore/DVI_TX/data/rgb2dvi.vp"
`timescale 100 ps/100 ps
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity",key_keyname="SYNP05_001",key_method="rsa"
`pragma protect key_block
U0dw3aYFMouH3CXEDfA6e/cdu9VXSxccK8hIIFERzi82ZqxoGn6nQL4D6R4O5q/+CErnyvQPKgb2
dATLwZUhnrhlzTJKbmvMljyK7GiaENbwstS1oql6oPHIQvCUyX6Ou3XRaG7ZGOfVRqNPvSrd8Yod
J5MOPRb7naSIietIk29pdfkDofyf7KK8Y1impOPHLYK2ug5Os3N++K4nifldA0kKXJfrGIO5tUwK
uaYKm3pHrKUGR72R2cAfEYSg9EJSSXKziyG+VVoYfagzj5tyqDQPlA9eXw24FUXZBu5qPN5C5i/C
xzrBIahP5ha0mqcHu37qwFuePWJNGYM8NgN9Ig==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin",key_keyname="GoWin001",key_method="rsa"
`pragma protect key_block
coQEjeeFBiYzfVU89oj5lF110E4FutGS+KE/zevm0VJsKRFp99UHVUK56DD7mJegkO/CZ/0xMfYX
OwtzYkiExdGVwHjtyucZpz7HyhyDrJIeLxhUZzo/6RN3axIztxHCmAab64CWC+tUrrgZ6UZZsYEJ
SqrRSJRLtikxqvRYv62hd+UApsl6YyY/NdUmhFrWzh+cA1xO3xKsITEcAg5E/cqiDmkP1BH3/0+F
m4TtYiiu4UxZDQdzz8Ey10T1hP9Y9qvl8uQD2baJF7aVFHTUFaRrqaz/XN+uuL6rm7TJcyoMzAEN
QazMw/gxVQN8++Q+nNsr4Oi9Ka3JtISK77fncw==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=59296)
`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
fC7HWzXWlOj3lIyq7jVYeY5PFx5QpdjytqRjX2ljkIqQwCADPnl0+ilx14F1AoSX3/l3qAWET5Vs
K3ErGGAd2Q3EMfKrb/G7PsdkixiBHoiU5sEkCQYuG5DbTzA9Xs9zsqr8AtEgHujydag1++m5cT9+
Odk86keVwn+oecJlMAS6OP3n/SDWpieX7gQ8jwuciXPvIpQJjdRf/w/9uVaMdai99YEh0jjLHpPT
hM5cNghxHleLKbdS3rXzG0Io8ddpuO8uaJ9E8RVTzcbAs0RVyElC3+FiuClOWEns+KE4KzK72Fql
eDdTIYvmIJ1WXtKJGBsCvS0QSTtQcnHama6wRUt28WE4NBkVrF1RIpV0ZGfqA7paQ0S5tQSXcmgw
K7FN0WsCdKPq9jqds9eL72ZNNhG2v4+YF/NLIzLTrka7uDK8dg84pMGZG+sEeaMzoq2rtAkN0JyE
JuGB0uzNYc+E1XlNQxSVIvKzTT6YTEbcR/6sER0oex8NjHuWodqhb0ufDm9D3/2ow8XZyxgpxOnv
1ye6k1KJDf2L09kiLgGW9HvZAYjhLb1QmNWRKFFnHiXa2yGnodlR/PAcoP6GG+RYG8qYe9BR82Tg
/HIvRRVa6KkKztna2C5dMCBp98SvecOp9BZxu6mSv5b/+gAKq/DQaWf+7XFCsEZrF/b5mIAI9dWL
+ZUGnG0elre3MHcgBljs+a6xNsdv/MTA7EIs4y4yHzgbICDjgKFGOGVSO/tl8JJnRAy1dilDKsKR
tuzew0zOYeheaE5W7cmOuKBhhcD5OaNyF7+eLC40ePx/fqT6mGD8W7J9zhCj4ZPxFzkQzuw+TFdz
2dU4cuzg1nOCZghZ4V64UQXa6bpE4decAy+Ks+tIYwaLhvMmmPLiGURYJB1nUXV9TtCk9bul/GL9
rC1klWdFkJJncXhyBx+ZhVs7uwq+zaUr4eFpCTueo74S8u/F2BrtHHRh64/3P534NIyxVbdfsu9C
EGy7ScwxxrQ5q+TRWBBAQqwpQqQuocsPml8LmL02BvmHctAj0f5wPobXVx53I57BBOdQOMM21W8I
gcFvgoLYWvwvheFBu7pAtaDPpo1QUYpc+fY/7spbWqnHqfC3++9gKCBszQ5pbLmYHRowPs+ujP/d
Z8K/tU9363wez3OL7IuMHGgV7vasWE+KbH8TSRStpKnWlKa0d6TyuAjqcfOGKM2W6jjcno5+4OfH
6fmsyJrA3UIMag2tSfd1EGMgwIT0whWeYm9X3zSfxNrQCMXliwcI+0fxDl2QgRICsBA5vt1tIffj
gSErR7EHWGEdIaxNn7sVHkuRc6oN1B4YNHBETRZcoCyTxsSzSmlcZpO5AqGgZZf/UltK6yxKSrEa
xEX5Cg1Vpww2CvnJLfkCB6MoTEZE//ndQ6lCflm9NPAQ/vUbJaOq9T+IyV90oYZeMNG17P+hafXt
vbgG00gt8f06tsCaR87ookQ243pMAavSTxXMjDMnp3gGfZuNNu0ZlsPWnWxHOB/EcS7eTOfd4z1g
Ed5rOQSiu9qWqekRUSDy7DFEAfUGOmbAuMudLTe90EHbBlXLdQlvkPl5RmMqnmeEyGIXBctufuL1
MwNAtMFAbuznzg8X+bDHyaXsqt38iKwKUsmHeFYjy0k873BQrkI32Ef/4eVGLfuK9dfkLRXhXdmV
amgxbpWXHC9nmPxmFcObXDCgh/hKuAhOnY0GcXID9HlanwnGIElfZja6p672QprQWLokfbgPXX4k
Df12BDX7tG57pgHzVJ3+GfHiu5B2j5hdblEzqGcIlv2G+asZ3KmfLSd+HYuC/ziIjziQy3Rxnfyr
ZPHA58zTqgGTip0VnbzOZV1m42m1aFCHEULTcp+PmLOX2jBiEDUTnROa3JHzu3kLVavtJZSFPdU/
J3aLSJXcYX3rBSb1GtYpjL4oCoawm4c/xD5yQPjeAM4YwaJpyAQJhscjBc6cmEFJCBRpI0zA+Tfy
C4GIVXT6MdauhSaaKCgkuwq5Vckf8fVRqukeRYwpEJXd4GRpqyioIo7TpzI0sYcHlwxyEy9TlmrA
rpgH94ZdANAKLI36D4Yw7ehOs5lF4efO8lmt/OwnnYx9QFhdeoCtYKQXUwgUwxua2cIgelz38MNi
i1+TT9IzOJQurYjCXyoXWOW9VDk+vTQf1V13UuZgOd7Z32QeUFuVSQHDn/gB+5VXnBQ6K7xULF+F
aOCIDxl4bmyiq0Ha1w+wK3XV9PAAoEiVwM8sICU6Z+u0LRQ5eyapKnmr/pBUqeWUFftE3nzsNSP9
Fu7RluZbSkDiXFH/uox8TtahAqWu/qlaAdbcYzSX3Y0ndzzloO2Xqj9cRyg/rCN+AQWCKEEh5Q+x
S+hG6bou0r//YqxE4Kr97s3WZJ9LygSp0yOqRL0v53EF/60w/os3PaRU0zILcs2ZaL37aUeAsy96
wPDWv7TJ0D5pNQMDzqjhcyhJ0ZVrAPkDf7qEC/aH6lm0KUivlsX9TEkxkrsHyxNzwz0DZ42pBB8e
WSatenLgLlEtgCB1oFoi871dpVRW0Wj1WQs8XihaO2Dyxx3THqlIj293Gi9qzPvATw/TzHbJqIBl
JkeztYJ2s2IEp6vgXSkiY64ckgRAAFdbajCebG0WJ1AOqYcJJGSXuCfpL4oZJUD89Nf/7uzQm+Q3
NlpjEudWRbE+0/hejSqV149hgIeGC8qR0LbE9qFHxh29wUhcnm85ttTkkMCgCNL1J5jmOdLC04xt
Nymgb2UNjTgIEjhooPAOn+UQMFBDiaH+69h+LYaLkGnlFdoUUYI+DURcFnL91YEjAw/W9tizM/vu
R5wSxs9OH5ocqCJJe4DI5aMSPz9ss1dTLBuggqXqHEg4jLtG/XnQlOhEGQQ6hZMB8v5LfmzI1S5J
xN/hBW/SOIVRoSdfFRzKvAuZgpVD2jRZpTLpp5i6aW3ozEfjmJ0YYnjIUvepAVZvzq2EciBjjRgj
oVE5h/ATSIn7pQkWHfnwcUxzTa1t2pyuxiY1p2l4BRHHw7Mve1tsSpnl2uV+EWawD5RHIkqSycAE
BZq5c7h0ldzPsBWxvOr4a49hAqU7iUYshc3jsZ8R1mZGH9GMNP+kdZNeArM/myQ+A3KnRJKznPN1
F8pbPRsY4+yLwLtHof3VOCM7QGVoq6JQgW8Y6RhmoJgJTujfY+SFu2eAdGGT97WY35cXNDssIGzd
jz5be3LJeYPIljVMZQvTbdfcqaP+3leMwRC0ChimuYqgrTiQPwfy8WVt6efscbC58u6KhSRCyKXz
rNece0S+XH+Rz1goNwxntYn4jK81o3p0u6qD77XqN/XJk/X/66/PzlnHI4WINYsiuAl2MH4rqlcm
zBOAvtTbR8ElL9VlR7El0VAJGrBo7RhpSgYGp8UueIzIn4N/fmzlyqLuesTVH/U5am26M04P8VQd
dYl2lEmCHzUeBxAZO+6tIyPsKiME3mtTuO1NEwRiuFlpaht5G9mBybRWVUhZSQYXaK6tMbvjjvV/
8+GkoolaLPzwN2CPzL9XVtU7woJ928irwK+dlqHvqFF+0ozYmjWCoUSeXFNrPDlcqrwx8Ghvtnhc
xqaBAF7u3fvzKulbwnOiA6x6Bkd8GeezA/SBTbt7RKilprPith9wIf7GZK/hGaonG5oIzP4hoJdh
NLR9SOn4anotlritksbdCMEDzhv0qna0M/XxfgsaNZ8mpWUsm4u+WXDjbxLB/8/q9g+iaRmrf1xk
1AmTkx+xS3CIjE2tsvd44aQhtK3MNDSLEljpoHZVD52wL8RWEU2tRVDcu6wSjG76QzU/kvNDe2lC
l0ct1F/W2VVIdYaC8WGKP2nWlb5nb4XSivKF0w1OwRv/h8j+/gVxTyDXKbb0kysfqXFRnps5H8U0
BuGK+eeEAjVg+hnCJJ0pRlcGPJsmVHjVBKff7ShjBo/tjcDoTDup/h/83KAzO87DOKkzzH6JMghy
0eG8a/BnSHQPNoJfLL9Lu3+dcGEFDJTwZGjVV4GMu8/ZfeGVfTyoSq2Rt01KwEXMJ5fOt+QL2cWB
RHG82U0iVb5RAhhfOHPYZcQm39W/ah5mBHV6E+0gcuVpMBZQJss2be/nPF+nMx0xzrOCAJjKQ6I2
pXHf6GrndZKLaE6H5zjtygRWA/b2duntoWEg+1Z41exz/rcKrXagNXge7N6ngBbE+mwh/OnfnfXy
TOZ++aRn+pL73Hxq0VRbLJgzTIzVyOAWa312GJ/XJ8qtSG0FbN563cZ+QFM1poXTe2m3Jkk3L2xD
bkp+IoWmE5iaaCT9l/HaHkfdtLGkz/rT++iXa23+G3qDQoRQ5J+G0UdyglP/HkQNg4zC33AnQUkZ
RvCR5raAUjmVFbIxKAxtg+jZahNQYt3+iORxz/fANl7WrpmS8EldXv3CssTY0Rw5eTPgKM+cdHjb
VQCse4XbFOYhQDZ6S5SucviO6xgJaKxt0fGpdseHnRUidaNHG1xsJ/WzPxVItexFzASEljBx2ARd
KUYAck9DYNLFjyPwak4Iad7wHPaUdT4UcGNWb6piNWguYpqygpD7HX9eE/Kh5pIWVoOuV6iHMOJ7
lXxMAyHOOplLfqdiek88AUqi5GsyNKiFabmkUl3zn0lAy9Ne9guNQBEOaluRhuuIZCbiVU8NZk1K
ErDAUpHRfRD40nHXpV9I+WXCBpTMps80R59gqKDQvaP0ZdKyQc5vVftFtVuWwedU3S2D5VkhZj5i
pHUpgNm1IoXbjvvh98lebAZPorZDYmZXp2ihSpYU/P5Wu4silePYvaaR0hPhwS2UO6BaAiyEdy0V
E90mHV4xJq2yzQ7kzPXDYBC4RFvhYhbym3RW05+HRYQ3PlDE4RzpYM/09hmDG877Um7ZI+eBBrmZ
OO0OjDrWV39VoxhXyuBCTqBS79p8XLTBkcvmtWVBMFJe6yvZLN7CCvu+O8OcoC2bAKjvAkLCScuL
arP/pZ9yVY+vdOK6W/luzu+IxPutf87ude6lMUKdErq7szNBJB8W7R0sAbHP30ihSKAYpqRGAM8B
Y9SaSGw+hUUhd7xX9UuHSpdy7YAw9eAMbykGr8ctBP7m/c2eRpvUDVtTzMMZHrgGgDvaCWpjEuOi
89XNW7Kur9UJHiGDe5z1LEJGcQmeclOSlNn9uRWOA1ZS1Gj563KGCyEF0XLO0veuYMPeuQdobbLW
NZrwdKeaHhrAKfJmCQFnxrAmK1dsUusOFhTrBPqSGxYcAdGp9uVEqyseYwvRTUcYpmApGw1zZ97B
EZzm3n77ziKhl8j2iU+FnPPFryOcFNLLlVrQE01rYpKCNcf14TAq41T4lZp/XbW6BQn1xZD7MTzj
ufxjR/sTu9YKBppw4TtWcBDZJawLOro4ktBTNamHQLKnEFRcjOfal5pJY6asE7S5kIsyqYed8LXB
qpvgJcY3nWfRzpKqF1HJd+qKn74+9pBdhKhtwbyyG+XHrhrv6GQwY13rwYfbUg9QforJ6VbIxU/z
Fb7YKNzNURzZXdX/quky+Bza4sIVOliWooxaKJjWZ/EAGRiFdlA1/ybjBbsjo7CXh0xxsWa3IVqm
cg3bFVUvkkx62czG8KMrrppwHIZDWKeIRAS85QOA70GNVU/Mbo6kYm6nXANBB/uFwtKh8xuY5eLZ
E0jhJ0Gzf/uXQ3vfmRs9bXcDhN/TCEyoR5owqWiGE3gxOwxOk0VEmkwe9HRvKfaQ+PLuVPoXh8ia
9b17VzYprUNfATLlqKRm6/h3/qylemjebshGymly7dJ2bP0y6XMmk2QNSekiCs85xAMIhStjtoZh
K3OZtmVVZ97tcYF8UlJ0oADxhlpZkugtjQQAUIUdw5g+lpSM9sx4IbnwqeoK+kI2a6tFHOsrWtRe
9sqm893aAwFHecoThoqSTD3n9a0H8ygWw02YTVJwDo7BT3laFBotJkK8KRhmsGkwtWUOkfI7hZEg
nfqBI2ycgrkR4k1bCSSZOwtpELsuVHeL05W6tl6MTJD522u4+BOfO1zjKsHhKogETUPO2Pbjsqt+
uYyKswRzDuO1BvaEREFiX4K7y9p2kaHLskUrzJMpH2u/LSfZHy3AEJXI8GRVayPYkjPycTZZ2u8x
zDM7y4/tIJv0yJ8nUFI2vPLb7lk8Uxf+uAb/Ml2baGHDWH9UKN3iHLTMEqw08rF+wEopk5VZ2WD4
vq14h9GF9aIGzEi7XRWnP5dU+cv/5keLCahYeE4jY+06kr4m4B5Tz64KPjLg2m1VSQNJ2+rsCD/9
zA/veXxR137BQylptjXWCZbpUN8C+dv85zkl92jrDbEW7R7/3OCtPYBF1LPlqIUH2b/TWQtSGoB1
YznyKnXzUcXIr3Sq1agvx7gUa8JPzUNFtY2ZHU0xGX3C/v2ZbdLLaQIZXWPEvYWt2TS7fhw/CnuQ
2PiSHpCje6b/ZRnYe1+zjtYz/nLCoyE9q5lNG1iNaI9sLNojWVrVamINV3uiubvwBjKtyM96mG2x
ncvDnR/I4FRccjjMluXH3ODWtYROyZWyTdrsPC+vGy7rNv3OvAhqjGEvQ1kKb+g+3aadXjMR3ASe
gyQoygBrHi2Q08E58l2PpqmgCnZQsfdn1lrqpHHcDaC6rMT2kdMGMOTYNmHy26e7PVcMaUeCHS4B
BxD3XXOG0MTbbqQsNztnbIOEdiV132FQrhHsDTgqMqBsN2RWaA4nE+6whkJ5hxbuPe1lSF9Pol8J
lD08z+ZDK9cxqIj+XoQnyLbGAZU/fBYuVddft2X9s6Ix63NBXSloARr5ClCLNYejuXuS4HXY76Q8
qfE2r5kLKzj5MLkzMot7hVgrURXyWgUzzcpvB9R8j3uR9RCDE/nnE1ZCbXICh6hC4I01JVFW2hd7
MmG6raWchJvb9/U8TDtOhq+R5TCUf8hSCB9mjFrz9t03p1YtiLB9xy9oxqrWyX1se+tzfeWHfMON
yPFK9Pv5M9sGSOoCtrSPMAkMrY6a6GT2SSr1ponx5DhcW9dZWwJFoaX+LcEWXX2diIle1VhGlc62
vM0vGG25sJJk3dewKfqUK+zGeyq8mnEL6PYkY0tpUAb3Gh4ma++Hd22oxcw7F8+IgIX6ZWZGV3EM
7gVK1yd/wsIf3Q0nqX2t1iSl7prwZpbQ9EdEsMZQMrbftYMl26AClxQ3F/U4U9eyHANgTsi3xu02
qE5IIfsYMUITlzGPy6Qg1VhoJNJvr0tYS9wutmoz4u/6XGcyJoBwttfFiKXwFxD12APVGhsxNYOo
9FDj9QX+aGMdF92sYaS2leIbqKv9i8CM0JPjmaW4+pR7a4c7MvCYBuyV3o0LliLAfxfAZ0Ya8vj2
oizugE2FgfmttQOYqwht3omwPFImWUckNzbRvN//3K24RqDlynpFEqCT0R+1XlyF4Kf+qDqQm+da
oBfFQRgjOSwc60S3gpDHjemWBZXvM196/PjC9aFI99a1jF1OKd/gOeYnudEqedMvdaI4YvhthN2h
EbC0TPA5DOSOnGwrmTFBH1SlhYoGp7KwnaRfEYhkZOJMjbH03zCAJnr9flcu1P7WkzGs8jjpg58C
0+3Cw6GmXe1CP+tXpe3rLRehjlzjYYHD3ox4EO7Su3Pe9cGNFUYacywr/Zty2n6NGF+Jje1blPeH
77OfwfDy13Uz/q9o6S98Zs7OMSdtiBjYWTTWI47TzD0Cl7pW8h1Nwl/9H/pobncLDtB4kY9N3/QR
ndCtSNbXygjxzyMvtfhaSLPV5h5P2G/wYhIGlWKo1vi+8sDC7qfZ12XfnPEqY6vI6Z5AB+qQwrGK
7uzypIW9DEyaW3TKExq3jVALDOsxfI3Y3U0zFCohYpy4QQVXEJP2pjUPed46fF+iNuOhEbD8iDHC
56bIDotziG+TLNlS8I1x8LmeB0y5IWn+HEKhEXnMn9FORx35r9EmPi63V/SkDtIJAMR6FIFKYxEH
YYyrlFSosmPMsIQuCXX71s58kG8gIANe5e9EGNZU4YX1AQHYBGNG1/kZeHzmj66Q5lXyMPxgAElb
5w1adydWZBY/JWPlttdV6+r5qmsm3wz8Zd8ejMApAym8UU30CoMNmYWNl8lqaUbIQPVxo8QnuI7i
svQf75XKEM2lF6uJSAk4HuEjDv9pW9udoUflgWpEAmfTTb6h0g7+V8zicLjRrLL2o4eSHyt0OVNX
RvuXHOj665CvJGU/3z37JJbooKuEZ7GPWhPO6yhvDmVLvOg6fUpLgVLfAmy0AYJVk39djwERg9Po
BOnex56dWNyhFPlcgq+LCoB1XnPa6vBDXu8xurJw9VTFZ1jy46fjXPSt33lP4hyFtgRuKz7qtFzI
oLyDvTB43A7BJUJhb/KYnUba95FdtWazOwH6dWjbTt7OO4ZO0f64sFH5U5lklOor+VJChQ/sdAMr
aJtQ1qIu7lrX7yDRAUXs7ORQQrBOVFBRrOfbHPv5i5joDKU1zYmRqBPZcuAkWD0wXqv7s+9/fzWA
Q7laTOBO8GOYdQt0dffGbkfuHxKCBdo56rF02dd/N1zP4Nl+ERNMJH38VGbsQrVMeAnJlXgSB8ly
H6BICcHnSQfMLW7Tpy/Qf9cutS+3gSyZCXG33ygQv6D56dFIzcYDgXOm9MRMWVCMe/GORjFptBhZ
zdqrPHXsg3cFGUWk5yMc8dfh4ofbYSWZ7XcNZDCAQQhh6zeEzigyGKcJKIoKjR5CnToXAm7azfwW
IwGli1E6W/YOarcoB8f1G6NOTRBxbTEP1tr6nXqJCP4E7o49SaeUhyCSVept/qDismggL0+HQsAs
vKEFAQuCquyHiCq0rE9q1St0t0EFrP7aFh44e5fZFiEF0IlrDtUG72ypuIweGADOmN3GecZMM918
2Q/tt9gFWXflabe4uVf6X8C6QJgrbsN1m8bxNGypb7M9avjvfUTLpR2SDE9K8+e+CzpZshfXXtUi
gbyHi4bmwEWbZWbiv76Fn6Dmaatae5P+XPic+zN4HJ6Ha9hiqqNziyRpApNVYAqywh3hTJZCwHpb
l+q1n+F+PvJvsHXkJCO1NtfwrrtH7r/Q532tfzDLmlRaMN2R0SyDA/OMvSfo7/WVXbnBobP9ODTC
BeNDk6/Yg3bzdTuVBdMd5HUqxjCUNpo8d1+nd1AbVgIMgBqyP5AoPNpfbxDw7U/5QIfq+ORLS+Ve
cr5pgjOkMsf0/0d0sHKyFRUKjpQwZ3dyyIy4mwE3AwaknJ6jBBnveqlGxwbo+FpYdEhLrk3NIsxZ
Yl/HrcLjmou3zrgWZwehqOwakxBYWAnSxERCbfthIq/PhsuXFX9S4pSQvs7KzZaUXPqtJFZ9vGVr
jKD1BjGe0iTilkMkark135NjhAPsQJg/gAVWCjLxSWCzgSJUjsvQsDj/1xD0WmzeHToBal5jrWUb
DxOmy0tEEBPpcN86fvND6ly+30zmHvjAmPn1WzpcTBZ0KK9cJDtr9vZpjV/bWpwWAsqtrfVUCVEx
FxHywlQmryQbMWBXgtcffcr9kck4A4kSFUSgMuLWLCx5Fg5tPojQ0Tve+ySZunawjdvf8gRIHnOI
YIJt2FhPVd6VlikrLsTrFm/B7O1+laJYGugCWP2BJxvmVaOSYcG0Gf5twncYipUxrvsX7wELTTDg
7u09DX4fk3n9sza3jb1g1F/LNk81tHulj/vc5GgBTB4/wyZjJ8lmuJdgxeRiw492Uz7ym7Sw8G5R
TBJumL69z/VddmyAq+o+j0v8NoIbCkl7uTS7dnkJcP/a6cPwRLgeIfwEJJEnx6s7DzwskIQh9je7
hjfhohD1Mh5ANFNAmnW9ZrGFnRqqrlemXE9mTXPd6DrriA1FSH1oGQ4BW2NeG3QF+FvOoS8ihPcK
9E7H6t7FBH1GRM0Lod5R/g/ifAP2AnVwkNw5cbJ9g5N8Xgd0hn9GWbORQ1z+XdqGJTDJgW8fj0pR
m2jGFk3yIEPh1HSz5xc/KLWZmAn2G2NG4vkXmXrm7FmIJ54Lh0wyV1KK5Bl4ow8oq6OuxS1TsbyT
FIxLFuz3LSbuWlf5nLr41JrW8HDZTs+DtjF4VyAN/FuJMBym7VNpbeO0m8GDflYZkB0PRK/m9gCV
7ZyT2iERLXStkg8EZwkD26SLreiDcIM6/gDB4S5mYVSEzc0tmiWqcaKbQv2Bi8JhUHN8ia6o/RCB
0dyGsdiyo3Tc75jp3nIvOB8fOwGbbl6qnWY+84qe+9kAa1h8nYV/mpnQd/7jvQanNVHZQx5VOslg
IkqgMgEHJexODVy8UpV0DmBbeWVJ4ABxK1Mc+xiAU9EMhLMmIOtPL4P5bj1wf+H5eeQIrCHGROaY
d6pjGOAIEq20qdAcElKwkSXeS5gvEvGgEhvLB9mOKxtY6VHhx307ODCjQKMlubpfiAuPQvaDfd8p
fyiXzpiZv/ll20GgFAhT68tep0tJMBXWER07n88iQCzAtA7nFzUrexmhEtXG6LSvGDo25Wda2XiI
aIExpBJsBX3WX7aSmRjZpwwJBckALZ637xAATWOIO5p4+6ITDothDe5WxzwAmybS/IEv5xjpogBB
bInVys06OUUia7dSSo1HKPUJp8sUaN8ckzSelUz3tyUtxMYJ6HcMyVdhtI7e7+t5EseiQjsLRAsx
ZWnGb9HVGvUO4NibjDPRnXzVcwv3Zq5UmsRIOPjWdSmqYoj4VA+VcuGVcmFhbTCwpx0CyzIp8TXs
+atpMK8jTXT2tHHVdYP4F9oittqNrs189tpD+hKRjegY/88QZKFdIL6l90qxRlyEK7n50KpY3bVz
rX+vZDnh22Ka1v3MXa1UGXivDWinYC4ATIz5bwPLV73OGVBXfh0rWFAfQzti0sEjMRDwPZgzUkiv
0hyt7yZRW9QRwP7Ig0etQR1Hr8+IYWL1Amewp76nTRheTxCvXI1UT/ZOzjUQkRtuo1b/HNRnnqXL
bX1aUprS8TnQDsG75ldKEmLxZs0iNAt6PTUQi4TlH/iqWiFtzefkSyIRm4f9rqkCgr40ufeI6Ufo
w6O1ITtisegxhNB2N6ENdZ9AyFP2zGkrO4oQvKhElWBHYwdRlNqhsErat5sG+cBH3Q80CgUuDY4S
hSqMy+U9eYcSr6ZLVnaSqPMoagEZO2GwUkYUeh0CHwP6rRHouVrG1SMGjY9g0f5MjUwc1wmVwnY5
RyXpDJXXYDElnGEf5CUT3ayL0roNtxPpjfPSQrcNYDECDK5SbBnbByP8fzq3YNz+zXZJk+tWLvFs
XRApq0Ps14wMLzZUevIOsIZ51mfEdh4KpuLtsVBexjP4sIlstXNd0z6yXpRMwV10vG7y8pteMuPS
Ld0AkdDl2GhCF4oEg7a5o7DPLTyoHxf8Re1WF2ozqLe6vAHj1hFX3fN1lkpM464ndikByOePXoL7
qo5GNro03UZCUvD6IBx350gOAodHWoAHWcWF6GB982J1rtUoFvs29M0E4Ul/Eyxs5NezzhAJXHGs
Xyp5ua9J17AVLKD/6t3VDykxoVrGTVRyofidnuIRBkBf7NH43n9kp4xOSPhyOCJuxz0bJ5aKMbmb
sBWkRFAqekaR9uQLLnbr7Gj80lndSewqHTI0cRPyKdjqzcFp4eF4yyZMcAFZ2UPkAYHauIAUGj3K
GLBn1HrQi5QeeTbAs2i8mk5VHvY6nxyuqqar0E68mkCqWLrb6xlKJm6vCaZfc2U9pdhfMkV7mqwD
AMB2sp2IgGRwgcKqqtCN/crMszDHsgkgDk0kttH3y4LBAAhjmuHGkUxV4IKKKkYx9rJRnJVTq2rt
j8q5v9C84Siurl8tqX4xtaIvckRc1SPKTGNYVR03ozhqSS/FtLO02OAjkQKdbJ59vffUrddFKA/K
KbTJNwji/gzaH8XFp8TnoZudzcRMTYRza7sCNvGDUvzvkcnBSuM8nn+cr+W/h0yPb04uyvNVnaep
BGVeEb8jCIFMYx+f+WyOqKk66LPaImCpyVvZE8U92Oe/AIKtL2xYlKgBhfY62uwup9wty2h86HtD
vLOl0pKhWBLD97e8ivBeJg0kBv9oOuXbc9znmP2YafTN2+SvSvtY0IvIrMHY9bQ0i4Q2b6d+K9Kc
mHeYkO76F1LIlm1P3ypIZQZapR8St9cAap783MQdKMV2fYmD2JDRDVBebQ2KzZzRKJ092q0g14kF
KU9b7jlRM290z8qz5q1T35OG2y0SQDqdBzipgmSBJO3XvjEtUY8pagC04Y4IFj1jlxOz8oFgY0BF
CovOAGN2w8qfUU8qMx09VlXp5+dbTBBJHhRETkUsDqB1fMKHFEcKFV6CssSteGkcKEdGWDPMZ1Nj
TuqarXNIZQJ701Rsp+bsBLVCzLFkr+3oPBVjpQzzom3HpOUa4XxVskIZvs9l8Zxo7tTs3cpxRB++
YXqm3R+5Wc6w2JmeRltskX0sOV2q4WyEhzwEJuljK+ZmJ4uCBQd0ls2fy2ug3WpWRGRpYtLPO7LG
U1xjUtIc3svkeK6Cn59+N9Qh5ol9Kzr0cNreMQ17Fg/Ac41NX0/D9pbwMTzqJF5zhw6reSWAHBHy
AjYpry5x3Wi7VzKMGhqCUswOV//ciY7WuqpAF7CNsQoheKH0LjnqTijLANVpIW6zygix6gbXMtZu
mTx8AnRwlNbVeSWlnZIiMK2UVdyNHUaLL94yFs+rtuOI8i41VlX9w+UEnoArVHTCFvrzikKQXSk+
LfGO1xe5kRqMFP1xTwdfmIoXdHv+oIwEzUd0aQL2Y4obYGjAtKIThPn5CTrMJJxxcqo2ldxWeENK
idSQEGKxcLVDmq4+kG08m5QgNcxQeoi+w8Em0G56/228UEMJTbkzvwgZA41Gfy3t69swFMJmwx7x
PnONMvlhxE4d/ypWUI7gRH5mU3FFRmEJRUedPSXQjBvqiyLzqii5SX1GdGk2/6jZ37EFuwF8iaos
LIds/NrlRMLpI4JduRW2GcRmMGi7alWyWVPPWJDIaKzLmoFFlv5T0hBBUImM7gYe0Hv4p5TvU87a
bfSjF/iycbiF/mQXRqzb1QasekulxUCbWYRl1rIBBIs0j5eFPJk+gCCbcE5fJi8oZV/xgKQ4LIgO
apxod3AuYnzCiFEt1wmM1Y9JXKg2Nf3rASSq5yp2GunItJa+9fC3EiCvo/8lNj/mT2jVdIZqhDh1
yS2EaLHD5EPD/HL6gvhQKS/SmnnrpiaQaiAhUHF3PlRGXvG7JUIY3bRebAaI2ra5vwzdFkHl98tl
Up0PSp8ZpTYs1yHq9+fF6sHOutIJ1037mkfeB3AXi5QX7cFUk7cOLbmB/ks2cnZ5RiyWAk567M5k
tO+dCnXBVNxUV/TfhfQg0mVTkqqzv6fTpDx5BR7kKy7jYskywXumhaTM+K4xAgsLei8PRKsgx+ox
XIMg4AL2SW04dp0/uLPm0M+NCa03NMZ4izdGQn0qv0LcOh1H+8+7ICIygEiYrk6f3EwQApnOQLiG
KxY96ZDqrHFCz+V3v6dQAD59UzcSBwDskz7gAoQAEk/oXDb/KrA8aZWd7EjnK3H2Bqhd7pZzYMTd
BUnGt6prk81hfFQJTmMlT1I1AUVQQd3Wdohnmyyb8TgWVrRReLLotf/XRQ0YMd6TPMcDeUDWxb/U
kMfy+a7Uxa+6QIm24eonwi+zQLKoEGAB/jab2VxQf29Md3Mf70V3vYoUuIEL9DA/OSDDfA72v5ih
xZKPb12VdYBqJQxhhZPjhD4M7VhEmNeVYGjrbMviwe95trxrd5SpGSeljtFEOBG1j0NQbmNzvmNR
EKD6L4UgKHa2LNOIO8eDjsG+tKo6ScofQg+xmK8Mtd5fx9GGpV6Zi7bSAUIMPvE7Sz7h82L1pv5S
/Xk+z1jF/gtXF+FFLF6inthduVZQBUc1Q0nXzfgYYV4qd3hIdG0jtKVy8UZxS7U9V5dV3/COkDzh
N9j/+4OaP38Se+For3YMb74wdkWHk8Fl4lVfDToGL6KcZ0n1Z8h74g1N7Pt2AsosYLMZOYCZ5TAs
GUCnkhhC2IQBkBhQZtY/B9UF2HMIEfmoR88PlN7DgKg2xB4ip5AKXJbFipgH+jbe0XB10P/QjqJO
n45WjfQwzHU8uEFJr6B6RHDs3hXaYGh2LVxJLGaqdLBgrISAeOwfBU8Ois8OsGai6U7qWTpAs3Bb
JwAhRvEsFQlW8gKO9qEQbrmsAqvgyszgG3Zqj3SgjPpYKA7Csw1EzY3Bzs36AQHUFXX6QfAoZMJh
CuPC9lR196rkNJiGngA4MOIFECCBdRu9uC1vdG9YFtpLA7ggyA4x+cvrJ6SUBJ1AXct5BhbWBtnE
cOOgSc2jQcDWqbtky3txHwLBcuepoV2dVl8nSe0g4GXc/TzaIFLANUwf9IQNx11cDkeVSKlZtEBv
gj83a8D7QUiS5/tqgROBW3gPqSjl9yP/053Vt7Hb7R7dhp0SAAxkSq5Ebx+PTNbtKvf70xpsIzMS
PhkLHIBVN7WSCdFaO9XN1nabaGZddfhU1DOQyB3ikeV/a16VTGKwf2yvOM/8FaRKOS/MHLteT4kw
ngPw9ncyIkFjwWkAJb2ZgG0fxZQ+QUzEWtpIlUYoP75hEGr6NmxxOuIzKy6mTFFAaktWkPR7JpbA
sLtrCS/47gq07POHPsIPGcs4vMj5nv3malN0kGUAG9ww/iB96VPFmfiUtrJGDp4y9SSeXw8eAf/C
ztHb2jTvE/iPXRFggUEZtKUCkMuiU8jaPwpQ6EdoCHj/TkMkxkXN3unuy/cg/n+MBjD+hhFVSn52
2CbsiAF0xaRNmWgS1KZkmOVjta0AjftH8mndJDABQl9cYNb3+orWGUaHyslmaHWoAxQPhpFv5vqh
Ac5bpIA1eAQkJ6sl3+kjaO/fB0/uS493aIYQMXb26/FHz1pdrJnp3nXZhW2FbwVGpo1mjYHWaunK
NYrl/TNwEh946YHerYrJ5BozQcnOLFz3YWI1v00djSy4nz+Q7l0/16DxfHtjWJMieaWH/VrrZBBv
a7ip0IcyQkr0Sqln+YR9BhohmXd8V6zdEyHd5+UiYFyfhb/Tl8P9JrC2cbxDKiiZ7JXS1WiJUapw
DzDkPch3XnIltXwpoVlwB9kkDuYQjLWoyiPwgTYCXf2a8uoXmcKSSwk16sf1z1EN/iS4yan6FsGu
CLB/Lxgjbiqg4A0jrzw4IrVn6JTNfGlTXPmI7lKai/AYREkJAsm/ITRVFo+Mg3GEbG0DFXE2Abl4
rVlHBTXAKaOuB5Ref6FDl37cVopLEoiQ28wPfnsCSPxaf+ECUmmHa7AWdFxnjwnB6gaVVwgBuNC5
hOofSj/EoQbdnR8GStatOrnzBTliqozJ5hp3ORjgVGzJLEa04r7k9uCw0uiIghi1aqmr0ZG3kXLd
OzQwDK7Tbs+FjckGSccVmYP8lAs0LIcXOh0mANmOaHEvjq/U76/ecjZSEcAzNyGQC9OFGc5+swTU
J51+hFOgENfgrO0ann3DG41i8N+fXRuVddjN0FZ63Pr3pBK38lLMtbJIbDTdX5HYHcsVt+18XRNw
CMC93FyOgdIKGZdMcLwgSPJcg1iFU5+tGIhV5k2qe0f3fvZnISNJ9XuYKZ+etdbbf7VeDoBqTrX7
0q54OnBUvp2gpofEbNKMTJMSW52Bgk0P10FWtG7LP8vZAdJvpoAefEi8DRLAUMP8GKpDRIG8h+RQ
bSL0gafmYGIesKtkcioKUXNL9Y3EHqvh/7/BhMuaVQVO6KgwrrojbHPp1sfdklraS6WvlrE+M3d/
EMTqUCpLgTtKETOXwPzBk5UoRZsEbFJH0MvR5Vav7rxwdCLq+/AJp7qhLbew8I/Lff+jD3yL1wO7
csHzHfMeiLUwuReH4G6igs+ZqNfULtj3hRS5ICJlmgXqulYoreUU3P+BEdjk4lx3BVeuBetqr3lX
ds0EurLkgQth+HbYxwxkudN+5xVE92S6y5XioWebm1A38qVtaWNP6H29gquHTgXuxlgB+LuOFP2V
KkK4ky1TYrI0CnJxDS4d+ruZQEkFaC88HlyqQks/4AHGDFdPWY2XYyktgMVD6uyPaEiX++nmfong
PdUzGSr5+22NBDNh0dfRIDnlery0OZ1UaIg+RRD83yyNm2s8MQSKQ9fU6n6c0qkE+6/ZK7hEPWjY
TX9We68AogF3LKAv8ikYwxb2TMQ0CFh1foDUTbs/hzbczzY9uqwzkT78k4UpdlOrDCW5xeCUnhYW
EQMdqFJZ4jcN1xLUY5XIEdbCofDPtgZJJXRWXwYejWQH9wXjU4WJJI9Q62SLv5m8P/S+0zYTSVhZ
pP8mAI4kiy4C6H29PY1QvR69Re805JB9HffKP2nyzKUK/ZGa+jMBCJZkSeqnSLzRuk7ZfJPn+lI1
xRcAwX5xyz/Y3MFG1MxNFAbDsXAhAz9UnN3bIgRIjSxJI6KvLyEJ2SdXfLiU42HFaGKjZN85tk5d
6Vjei6W9Iyvqpmhucrv+L6AZXpniFMJMwrSRFWTEdBhvM03monK1wcpCSxL6y3R9LDjSZ+z0scx5
MHy2FK4EsNPZb6VSDCMrP1iTgakVMLLXBSeSMb8SXSRbfMfqKF1+Zk12rJREq/3vmz3WgH0fXRhf
ogo3Z50+OL2qWWFjODhF2x4pDS84T+GmTAJYVF3bFOs2QuahSdQ7Zx++LjlYWlTQAmLEntO0C5tB
7y0zieeIIbxCyPZt9yNL45l4S4T5Ef020CC9BDWZ4wdtVtIMFtXhqHElVd1wovDKvdqrLggY3mGH
ng18LTX0Ikm8EAgUP7UdLwIg0K0MbeV8rnpVBcm73nRYtf7yhyZaoERnvIXyTVGm2VVDgf1yiurm
fT3thpa6wXqwycfmpDdg8IUG1nF/2EfyodJosAnmPOxiDGBH0hjZMn/qyUUs9ODX2ridhNtKyrX/
fUpeII7uSHptpWNnx+PnR691QFPsqhUw2x359ze44OfbnYxtpDohYNGIHRO8dnm3Y4K4IWPg3V42
uyR4fQypXY5gPrUX+bxGD2zdee6sn9tw6u8auJ2DwusDIG1F5VtjUabnHgRFenCbehH+xgDiwyhJ
Px4R8UAIHvuKfDnL1Q54G9fjlVfkJRr9CszOdMKstFvfRNwX1iPxsePSWr4ZwLRN7Vx33q1SNCUH
7sVIOEJzNjWKPlGYFkj6LgEVCKEndxQ6IHbAxqv63nl5j8NQfi5q+YPlz0x3M9/HhQ9wJvXdEizc
RVOQMrimzaFY+zOv7b0544pBXrKAMxmHM8Mzle+NTDgti8WmtXthHnIvPidqwZLFE0/NoC6jfcOq
IuYOu2D7nwkS/QlsY2qu6O8qpyQJ5JQBO7RQAjYFm/IwXoW6QTC1A1SgzeuYGzaByjF+a6hgGV+H
es4XyqluoNeI+CUE9X3la9v9+RaRcsnz6ZIAdY8NbvFLWJdzuhYa4ABPxKywNNNVOsN+NDmvkodi
H7122F38GUt2jJmjZ6TwVNR1zw5y7VHdyOXBwUThS2Ohs3ARYrqv0j5tCWRymU4FOWzfc6gOyBQ4
TTN4jDnsnMimYdlbjvp9EGS8+PiLVx5IpplTpI9o/pNELxL0s1Phx9nOad2BNbF4iJFWr5iFtFf2
LKCoBiwew6xKH1A9PnStwA0UZdyj3daGe3tk//c9kWmR07OiO2v/qzTJ/JJUyoj7gNYIjK7tIqWq
57dcQ2TeMzL2M7F1SqXVF29OMitZV6pcBOnDxHLHB98dk/st1kVb9394dZ2hKvQFAksLGIyJwYsk
R2nebgIMpt3+dVIxRIF8Q2AjnBDK8u+9mO6m1Evnvc8ln0aYDHtbK3yVQj4ylIL59i9857oOUU5E
Gl9HNTOiYMcnwKK/bRgNgeDnjjv3RLQmhL1RkFUGZAIaDUpMwBgiVP/W2oEjPk7Af9TCVGWjcp/U
OYJrGtgTb34P9iDf6s4kqIKp/6NORM1qRrsTE/GcZJKQ7NqQevijAXoKxAMlRCGQdyG9nwSm07qA
5kakUzONj7rtPRySeWvU3xfije6r41KaxKbZO5XpMrrkpuMIp3woBVA7JVlEsJvEgcQYHbz4e5u2
QcfnJQg6WMzcvjFCP5wf/+WGsx5LrKP4DKGdHNCF9xswhp0vaa1t6A2qJd6gZ+TzIIC1L3eQO2ib
pUkkRXrIZ17TlNmHbrJXujzrhAlZUoIe4E4Y1KR31kQVYqGsVgkOhu8QTYD2g+5NJNUOrt6q7Qmm
fDbYoD8Ag8mXBIXExKjee6xb5AQ5UdqiAfLjq+0/pVOBe/yv7KBK4woqhz1vNtqycJ+fD3U2QRYr
RSIWDUk6FKY9Wz27QXor2M/wzTw+pWGMEDqqjO2Gfr1kPrBK++ZUIbHQ95Flh/+QPxIRbyRQfokp
vMn5b57yId3NgFGYUkoCF2LedvRZ+cf8/yz2hpWw858NlHSmExy9fqLIL78coCOb4141/rdqSui0
cXpqZ9Hkp7LIuYGVisl2UKdAedUnaCGmk3KoU9VtNbndtKzAsC8NulRTszXqTLt/tn4+ZXqVS2CZ
B+vIbye0FcHvPdMbD2mlJWP9S9cCRYbxix70giD1n9nTNFxxTvDBo8eRS8kWd6Frzl9Ml8qzOXSR
MgurE+7D9Ztt1gUd+dEJXpR6pVwmXC7T8h9ht0tk+eNJxxAGFi5wxoLPFPC0tWxH6GwE7+YrBGJ9
n9GtVegBxYfVlrNXll+hLD304JzjyBTkC7xVGEwtc3Opyo4gBnVS7rejeAEylqeHDtu3R7S2iUwH
3H0SqkXnSZ6eeZQgo1j/gKIDcGYTeqVPwrjS5KU3zQx67lMhgTcx9wt64d/igUyKnh7YB6z0g2FE
6M2LpS01zz1bbM81Eo0MSS6AQnwTta2NZDY0zjGLKzWlX/K0iT3RLh9fQvnJwMBioMcbtEX5VOwG
wK9dp6VxvTh52EoQRckDEv6E4qWZWP89nqBMoTK9YxrTz6thcs2nlnesQSIc3eQVk0vfHJ0DCVUr
SbBwTU9+hKgkQ7u7zqYxbjVIxCnkZ53lzd8eORAL19f/P5jJMskb5z/rvMFXZRB25B8tb7P8eKEd
UirwcCxY0qiYNL9YsfYF+Sfv1doYV2EmH7Pcm7hpHnJeE8cNTf28rjhZiStJHKcJLAhPteIBPmKW
q5UagDFWaZng/OxsRt+1wDcFASUHEJgyDWxsJ3PZEBrbxKAUAE4lIqBpe49cdD6G+RaCbPUMJUgE
GN6ngiTS0wPcEMo790njz7C09yWIRFDlgY5FLuNmbn9B9DF+fmRQjY7Kz6TwwHWl1ZohKlscMDTj
Gi4Avw/rs2TNfEgj5+5cZPKprSNacY8cbRRd9QLdKSgMQMJFzpdSAsxvRqz+wlzVwrHmPl2ZWOXo
8r+nbkk8sJeviaw0bopLrVQ3blWJOVkIAUfewr/EEN/PbtzpWkCGGGAEByA91vvoDzfd5eA8ENm/
I1LOsnSkr1m2+czsusxQfudu6UaiNPMArviCxxB8phMvV6vvk99k8KbR12xGyHmezBX1O70UYood
hNSXSOFSO8YRBxl4mhP1RZC3rCm9jH0evaV5/Tb+OhisrzJ97gJIePNizV3DpSO4p2XePZBkBA+d
b6IFuMci7HggWkYgACK8ORTI4fQZ+6GFvZ+Di+78Psn7xr3hxbnYXHhHG6mG0ZYcNy4Pwd0sjckg
YDZRIGkNkTpchc6OQLzJM+7tTbJ/rrDE4py0lJZeyiGzhO5c+9gKfEktC+Lx81h8HH+u1XxKjk+J
Qep+XkG+VGJ5OYnc9LeYXVRLu2fzoSAI2QMGkXYWhOlFa3bITqZ9SxW9r/ICV73E5zGz+OQ1ZgzD
02rfEYLlwtnb4CLesnFXTdUSAah3xNL1pauouUUxDLkOjc3r6QaqHQl/mMNmHuOX3ZHqXUwcBsT8
Si7JMFCMFZaI8ab0z3gUcU9JPy9V4KKd5Jl8EaB3Wfu/k7C8jZM+MsbwyoqbfLTgNwkTxcAPyYF/
LpayAolYwZmZJZLfb+T1Tp+41PJ0N8EemqufrwS3esf8IitvCRT+XTTgaT6+CoG+H2DH5LiYDsXk
ll1Nu8NRqFwkoirZ/P7af2KZor8pva7iEJN+L4DEK6ivWRIuqYGAvvAlmrzWO8ezKu1PNAzcoo5I
EycxjYHxup5p7symqcjN80vut5RZioUo2dz0PXXy9hwAob6DRfOvPSujnL9P9+95xOJL2h+XpzDx
XUiz1j4YLu9H8nLTKUY6bKftlkslc4OZj1OEbnXNBUQilzJ6H9mJzLoCsRtMppZAD//uxTdpH4bF
kKI34YJI852RuzgzUf4+/vndVumfrBpCmD9UsXC/w+JzZPyWH/m638SRqm46oeq5+a4CH2wwlOp1
CpU0gVI/KY72rwCQ98hmT9QGW5YT8H5CBMgG2EUhSn28Iwn8WS3Qg8mLahronSq0CxMQZsCvn5Cn
CfN9yVBdpMxX01sqnteXISmOfJWhJO5AM8vtZAhshPHCcJX1SvX57cJD9/YegmXiRv99hGxvHs7o
fGhLTbBe/Sqjwl9MeJ8qARlMlLC9S7cGv6es1hFiHtvXh26ELqBv5ztqCKYefurgMyMm3iWQTxgy
WA67vJZBmg6w4520QLiXbdgndm3hiWmh0hx+Zuv0sGs0X3h2+CpQq7h4dk3+OKvjQ7W6PAelvfHl
TTH/dTPjcXDhEvWIu3fX8bqC8XmnoJf8eyULEOafqDgdExcjyKvAbwJ9d9C1lyzwSZPwpJTy5w7H
LSUGo4JL6HUs8L6aSM7owep2yR4LqPrkd7whj18dsBpGe3dVMvPUbc+Ady7qqz56K2bd8ezSVVse
PX5AHeY7QtryRuQ4QtfIirLnA9drsHBC1nOKNfletZPWrDapxaAOyFLlchvDYx+gAYjDyZciIdlX
VhtWfJS9iVtYGYy6VwLf7ZH1R/sGNElUorNwC/cmHc8PpiTi9YbMpHtT639qUIul+7rG2mM2aPPF
BaWHRrGXC03wC/KxwkUgCVKbYlnQH2z33rAqiZotc1d9UteqzuYjbMpEV/UbPWiS5hqxy8uJ8zOR
Yke8Y3BC3XzufLsESkSQnSSqAD9UfliT9U4MbK36qKGSToyY5sXckHXJVCfHMjD8N+XxMntFm2Mj
lTtzM1E985U3A/gSBBrr9viD+ab67pWbjtOcP6nylvzL5vxyLYbgzoZrdnQeW4QkEy4PAMyd6ENO
U2FeSvw0te4KM+vDyqHg00d2DVWVQK6F2Fl2PSmelHRuXDueXi8+Mdq7psvv7MDZovJ2AFy6y9m9
aPM2XEUWs9/BNCcJweJhQA5bdOdwr5qUKDM8cTrtN5XAdV0NM6HIl7X7I7/j09GEem3vEaJxT13E
hnqce3jT0fWubFgrTP3cfKw4XIBQA3O9zp2xxWI74gjXdE8jmZIRLRT9duibsi0pJDLw2iwtCk9i
Uvh6RSTGZaaCEyd7A9fh5Ezcq//d7Yw9sGo7qPVriSfk2l479fchds7E7GnCiACxQTFqY00P1mto
1XuzXfpVSr5OVjJmeY+t4kwAsvL/n2Dt84GbO0DWhK6qixzoPRVECCzNWbe4ssCRRt35mS3R2MWJ
18Z99cc85f0GEwbnXpeRoeL1fJjc6BjgZk2RwwBKTeBbkFS7C7PHbkEEPsUDsnwhP7SCrfpSYbNb
fwHXXvmiZAButZwEfY7pDaRWxBCcHVQlkzhRNmG9dsaWSbVK03msrfvkU7QpTIdWy5qkQXb9oGhd
J9JaBTX7Qvn21KIaZjAhDmESswRLTk5ozJOidP7C0Q/SdPH0+PrPGWrZ9QFwv/32doNMbLqGsVgS
VGGIaVsuFZkPVfRztBE/ZZpfwf8QBrPvxzgZwgF1/gMBgTttWgp3vxFjws3lY6RR3nZwkUs4z+0M
MOQ6Tpx55/Hlifg131UGAM2A2y1/GxAqjtYtuAjQA7FYb5Es2oQpyvUI3XrcGQv692ElLIC2M9WR
47r8M6NJBmdbH10yhU/pDrEEVt4O+PVJEhzTVWudxyQarWiaJEGypP8+yv5vgpNTeIUYmTCzZhvz
yP5rwifPyaUd3l/nyCS73vbesxezAKf/56HevzeTO4Wy8E0+HLMXrCRrurg6drArgXJGppUecjYq
q1p2ZvD+sN9GDYy4szarHI++Wz/qcggKHaYFWEC+iZwy0IIJ8zHvqhTFaNDpAN7lDLOgoDSjGxE2
gFL5g+V1wAgvNICcrfVV50B//ZC38jU33LbHOyihu5uDoVWw7QbH2qFIv5j83qYgDDL5qPOup0PJ
ZtQLLNovj3bHnU4PmVQ2RkNKDi+7iuAwF04xDREaUIe98kdrYLWndihF+UdowKePL/ABUG+E89pL
W0U4T+fb2d5G3aPNE2jJhjOw8m183ArZW/jN2G6lMfs2Ww6vivm3a2kPOeHLBBivxKg9AKWIRkvo
D3ARdfVt2YoW+ed/7oOckfqxH3tOR4xZbisTuklzUsjLF5fr+j2+q4w/vbnTW/CSCo0MxUxwZmXk
f4r/Mo8fWTYeQH/9yGihfZF02cGvzUimOWeO3XzCnkVqna75MOgZtDWzovnBEEGb4viEdtZKwdo/
+4Ys96Y47T3oGWkFk1WEj2nvJ8VXEcd8RAoEcdYGSlsffI6aVIeO16m2o02828UsMzFgeD8n6E73
4lZxmdkgFcvtyLg8sL7yB5Yq0xV4xbkv8XuNxJOvL4t77uJ9wYafydffouwDO0Sf+oa+kbQo/GxF
o+K0Sa8elTDjwCX+nbb8LAd+OYhKCrCUznKMs3PS+RC9dT7udYwfZiA5FGYYljiTcFFdHjiwp67l
j0MSG3HPyKcd7cpm5csWzP3T69bKJAU2hKyeFJM1wDmhHNqY0hQMYer6IRenKGiz7DR1b1VyY9g5
Ez2yInwcBNYb4ZGSuwZCMDDnRKIf5T6FL1PfDEFyZejApjoaWJ7WLKX4v9Q23ZkTwRR7AmnomUVm
CoLr8ikzH38azJH6bDgvVjCaNl6BQ+f5PJCRNeT8RoWygJOr4VDb2SNpgv68aHNzVAMZYIeX3BaV
nw7aSTcUg0OhHJbzLruNLr7bN1dm633qC1n6HJELQ62Yd+oIZsgtUa7IH83u5gAqtG9r0bUOM2X8
f9A2Qic8dN+g02qwOnv91dwU9tIaKWysVIBOVFYGPJx8sHlFnSF+WQ4ENK5PbNu3ubyVtt6bu9z9
LBTeQd4k0NyAsvVUmsB4fABTLNnNUPOxJV2l0Ed7DqBQsCZQvWD51VwDEOoPJxasGzGLr9+tIr+C
X4oHNTiFylmXLcPSqU99pOk5K62YRZpfbl3hUZVCVvmcV3Q5GnpVt+a3qLbSByvTfXK7bBzQmuEB
bRVozh+TiVM485w0Zcb8plVoi/H7ol0dx4qAhEEYZ/29LgalYdT4ki5PMEMqLQkOsMfbzQ8AaTyz
1vfPs/wOaZvaeoI2Op1Ps+Ac7QZLUHYtq2sOi1V0HOqi0sri2yihgXqK0TKgdVcb+JH/HiwAHIQL
Sh2H/UQFJAaY3p9XdXSAUsvy37rc6TSUj6LZeU8SkA4W1b3/JBXONauB1ryTY6R1ZyAhdimK4NFQ
K+Y4SH5khyUhxq++MBowntlSD74pOHVSBRqz2t4Dg8bOBebHe4+13CvfSC+0bLRo7QxFSODZIi2t
CkMORcv2FV1EJJQe0uB94NVtxie3CIOhsnQE5a4UUvEvBTx13i4N0Toc0ToV5+bg9CCnoXqX4tDj
/aG+czQB/hgwBj0SFnYl/QVYquqiuIcK2lcTKKTVuES5rSOWQahbNcUxDzAGF7HWC9NFL+20sAM3
gHL1kjuBoJzVEFwb/Q8Ghjdy1tIpH6cUqCB4rpCGSFGzq+yKYhlpdh8imtU8myeL5myzRkQrugwW
JCcvCfDtaD+BkUxI05BW3av9riQ6EMZ9p1e6Lc9gLhwBHO9hF2utK/PeJ5y4LgYR7ixPbDt8LXs6
gWjVj3mWPt/Q3il0woOG+0gABsxQTV3sJLXm/0OSG3cb9uJnpLOprq/qtqGkFvGSONqTVk3GVsR7
5znGNX3gBl/yLzwHqw+yuN/uYY8N+Ntuubl5wiOzGrjSLX40NFpTfd0rQbQpr5MlNK34hHpOVntH
wtiYrJI5AvYsIih1KrR73UL1Y3qDgEkveowuIlgDbgHiYWFuF1QmT6W52jRzu8AjTLR3jOIFAHF+
hSUCIt12PZwCRjEZjNq0TPS7D9ZacTvzawRTXMT1KriQ+YpTku3XHP4VWySwz1BtttaxbOabsp1I
yNWgm1mD7quMJa6BssrqYns3iuYsaMK1PUrlF1g25aH3jZfCyyscx0lo4q129OdF4WPhBP0mp8z3
0jEDyY1DvmDxRV7xC8hdQ/XBY2MOtqplDj7Oni+/VmHwfMenVZKf8UImq7/68kR8mLY8m1It3N9F
ds5lHsgDdL7hhpNhSXyvtrfoSMeteaCI0ikIgdEWBXBvGHOm4GH+wZmbp7VbrFUjtv0zp28L/9LI
Ps6KD6Pep6ezEU03nI4wTylOptEJdIdyaMDy9VQbDbkGU1wGxOsS9UZFd7Bf6AsvrW5DX/K6Dhh1
Ch5g/LOZ9+dT+4dO2+AjBD6NLO7k1JgNnwZ4cLXJDauGlepPeQ8O2IdloP6u4JutpBjlRbtQ4tq0
1S56z/dRv1BK10fXfN1/TmAAqoz/EeVUIip64pjfO9cDI5076+M4buKyKyDFaPtoHGxuLp3UmyTZ
OQKhXyU7Y+O3S3lCRdZH3kBx6KxlJi2CqlIkLKYhdRDz7oE9SU/w0MGLSH5HR6GTtQ4VbZryO1oX
/1/QU1YhcA8Y9qKp4Un3Mte020MGowl7CmrcEDwmjmRbQFk8PaC5Z6OsPZ4wBPSbau1GwvFWBMeS
diE04yz01VOyUmyjzIHFq70fwIc96pLQXyzapD8qvuzcOeLwd9cVk+qlriKaYre7F+rwj5e0h0Ga
iKrFy+wvLhrWVWuMedK1hqoL33MblYrhy2hUp14JxUXsaK+JuNvUl4ULLlS1SGG3xU6c9kIStT3g
N/J+UlkNWbHDlkMy34ziaVde12HfP3V/kvVW92O+L+zDrAuVGmy5B0WsZkiuGYwsmX6+19uPDgQ2
AzYBXEXAr2G9C2u+mCzBfKr/7rJvPNHjqP1U/Tz63QJizarvO+IYko6jCmqIGBQvhJ0C6ZaTESlC
nZYQc4qvuX6iLFpugkMKtFky0e1+onN13HfoUVe/Mhl5ylSA1k3mEzsqAEwDmtzdmh9TygqHV59u
KjN7mjdtPP4HD+9X6TiZwaEKzvlaErSF8PAY0sEiTITEVcLophap/v8yOTZvQRb4DXjyRVV63RKM
bi9Mcfe6+JOup/2Fz8FR2ZI7YZaQNtUm8b30S2Kguze42VT7usgbiZpCCuTJQgrLX7odkq+1Shnv
haA1llGFlIpBQRdmbnE4UpfYx6qYS0XBzBVHu1slPbJITRuufVz+o/MpSiEwaCmjvbWxypBq2twv
eFmUp8QqAFbuU0vcJ3Oszcxm/xByCigukfX0bsjfRbLWSBbwdiXefEX82Q5YeZOW7A7OJhuQqcPA
khfmWjE9h9hKI8sX10H+tcS9CKEtmAJDPu31SQ3nQXDW/75JZgWd0a3kedZsbh/MsE1j4GSlNUOR
5yFCC015H+LaiHN2jIp+YWv5MRAIu6VNCr7cTjCwVq7GhUnT1boDqFAmneIwIESkRsnpHhKJMvK5
6wtCWMH2EG8xrdX8jrbzS3UOtQD3y5gmCF/qRylp0PXPunwzCjAfJcHu0Hqg8+euVagXxNEOhspB
UpI0LGyCVStm02SmVhRytgXUfZ02oJndq/bul1hxodUtUQPapZ0TN6GlTdO/qZ3ner40oGRrrZmQ
BbAk+CBBPaay+ftLFmUJPO+c4pQJkV3gaUKjGgleHf3z+our/S3zHSDK1HaiLi7+dUabFAc+/qmW
iuDPTpDWy0Fgb8d9ACY+HC9K54cj3lNmLXBSpTfgUxLMOPcwsx85t5GsJmXLAPhVDnJPFy3/IrKm
9nx62ziN3vz7KYQnYb2UTxLzO41e9guw9XUVE60/DGhuwdBhoYcI5sjRuwG0VIQBakcOFrYtJxp7
JCKZhHcrGILI93OdulVlSeyCj7ORSfDbrrIitw/bozJ61dkIuk8Ru4m5ZnKsyR2Kk9HasC7g/f8I
82TwhqweK1vb9Bnv40bgz12qNtAZTX9jHi0RU1Yl1fD2pUVDOGczJ2UcW2q9Ej6ZNk1lEicHul4g
lpt8hq5V2nz5jNpPLQftQeW6Se88FBXJ2jSRZw558EUav9rwhUxkpKdakEBNUWYW7ifFp7wAbWCG
JEKBuicAjY27bW+O5XOOVp45i689ihsegJlWXhtmlbEVn08ZDGZekstwOE1xhqYrPgTbh80OHKk3
PAAORaJ0imXX4YycihxJL1/tOrxD9239b4brVhfERumMe/2tyLDa3o51Mux4svE0aWanUnkuH3xw
qgH84yOM0xVG8Dsx8pctGINpm6HnWD9/ih8Ajcd4EvBuvgNGAihxQfO1dyEgcC2+KpBVICwcj+1X
Rn9U/RNMJwg0aIS7S6UZxEIsgNILxaxm80xAAg1mKr48DHsHv+7qm/A5bhlQzELv+Shke+VoETiV
pG3IcCR/9Jg/6xYCCK/ScLaTV6DDGcZh0DrXecNnyegZVfAFlaTZGI0BX7lOFHeoU0moL2hggNs2
ywcbc/iFfXckmBCr6koQZ5rNSZoHAY1311u01IZ9qpzQaKLfABLxqOGsGL/FoaREahlJBnDiu9w+
LFB1lvGtP0oAnxmYhQ0K3MzQK4089A6l3YZyc4SrNO570DbaFvOy1ogRim4SGpVk0N621pyozPfC
d/96vRszQh2P9IqEslwB3cjkYudFBwlKuLnFlB4UmS9kUtnMqAfAmJr+p1HmI7pDaZEey4/TSiwR
ezeqdHa+AvWfQaM2j+C3cFnqZz5DEUvPxXgL+uOhkNWPH6+aMmp3TCIVmDj2l/857N4PtwHI1/68
aJtXNZwzGpzsrwgqu6fkumf8/L72Z8TfEBQsly3Oyx7XnU5FdY4a2W27nghrlBD7nujmclzJgUE9
2WpVecsEFuOfVknqcx1xsT59ur4w/zKz48YH6i/PJj4YhPgpdk9tf+0tHk90iN3rphvJ95tX6T1h
uXq0gp/9wEudwWOk4JJJqGR1mNCGUVvzMNsW4k78MpB5kaiKTflEmumnoWNMQiG/UfCIiTSXboS5
fxTNzbrOTLJlaMIZxqFy0dW+msCx8a3CVyTQNQQ4QPjfJPvNM0ckIxJgJ9oSDMEdtHubwKq+KbZz
mB+KcjmA0lY2xhBF45CBPYvgt2fKzyuu3PB+3nPKpq70qyy9dAsimvvzot9/i2FXXfgz5vOE2v8I
cf7hwYC63FVHU0qDxB1Wl+lDIF3eEbpkCV+JkBGhJEq6s0hycIt+dKAPCOTHlJrYLy6vfnUo52I4
PlCj47pfJWrO1kaJtB4sCjANeNlDInd6icl2T2Fk4HzaYBP91A499g83DQmlwxgs2Usx2MfNUGbr
0VrTGu/Yue7/TMmKQ0HkySXIqBRwE6ogxoUQryDnc+U1CkGsXpMaUVhk+f8a+25+3CKgi28ENoD5
Xn+I3dznjka98J5EV6a8vx+GB/oO2klS0CdsxT0aF//tmUfEUIybGtBJo5lznhlmXOmDoF+plTsD
cEwVh4Rr5qnTyhBwEF0NaWm94rshlgjspbdEdWCF6CjzeAVdl93BKXmFOunG3cgrBkCh7mDk4T9t
nPbGjxznQIdfA6+W87uqf77C/EJTOqAPV8JeTFjEHDyHa4ABi0Gy6drSX2TIkmN6+09m92Nk2/na
7zdQWfxvHHP4woOcTVCBO3Pb1w+LgES4yXx55EuYU//VHfLeTAA1/yAATAylRE2u8M0meOB9oPUm
jId15UC8NT4igiq00QOo8SS2O4eHI4UMauLc+azViLDJbkoOT7wr0BYBCI3SzP/FHPJa/dQTYI6L
U3R6EmQO3kCqKpFrrQ8OkVBKuT8UFmgbp/lG8iBeO2JmgzZCfUUONw8ffEfkKn8doPDja1UERtos
jZd98Mhi3qDHshL6bIfmRo0mfaWel4bzYPgBbBy6LsjJGd+1ivehm3+mtK0GKP+o8QVvdA/csijn
CXNnTBlAqRJjTP2fF9o3wWi7orelo7x95vNlLa1Na1jHCGPTZTjIIIWZMYe4K4tswxGShVACt6bq
SvhZDfoxq3p0xwatHz2/6PV40OwBtadzItQ/b2cg9Ejsz7H6f2NHbGA71tH6Sl7LawxiIfMDCWvd
CXn2NoeVUWLV+PsaYJRvI/yULqqwtiZqNgkEOI8X4HEL9viN5Ug1XRj+hN+BrFbEwGcEKCUEiK8k
z/AAwsoh1UfSF4q7XVpLsgqB2m10l5gri+4mxvFw137TWTL9p0K2ndrsKxzQwPxs1z8LZdfrw0/Y
0wIGfWkpEAZAqwG+XZHMHWeSW8xw+lus2+bu2cTgb4iUMtPDZXtyPbegiw3VSkrz4b6XRApHrdbw
lP4oUZNjY/nJ4Ut9033APWzWm8xNVELkb1a8CFMpwxHugWZpqRhYutTqTfeaCLVAbqosYydwH4Of
Dg23rz6M7lV/K+MZEphPMgcnaOd3W4zbnhM6qc0I86ALYaT+wFIptxGRwCUHcJ8mQWDCAqAfe8kC
oyj043Lb5hoVcjfu2ZPF2W+/alYCktO/Cx/6fdh2T1PJp6ZlcMQr3Z/tlZPuyw091mgPZEfb3ySl
vSgXqT1pMjc6WP/BOnBEpEjv/81DuDdEmwmF7GeOPLgNqKqd1XGxpNhcZW0IxyGt+eEVBhvi392G
41yKcSo6O2DXr0rzh044iQrd6FnBaf133ZmZRbVUhGdZqk862rIJdXsgzqbMK4qZTePuG1nCRHXB
kTJEDY5pui9wWYCEDt4wJqoC6HYFOob0n29lltNvu1Nz58UrGoEqEapeAiatWFcn9ECSejwUcz+4
PyVd7r+z7xFQ2MUMuajrnPChq/JhHE+tYYaiBWWOOAqyabkyDEBKbrHmstlapWkC/C8PosR2DcKE
tJcpIs4zYbYpau+dax4X/aKUrPRjxWT3zBEoY08ZbL8W0kBoIK4UUYjVeQcsg28l0zpfwYpZVlTo
Qb2riPNiPDuroVvB9A6dJTzS2VfcJJJN9TAPIv6RT6TLu72toET2DJsLL3PGGTfrFYtI7oehwYKL
KZBHeRGVGTxxSaFHUd5t6yHcavU2B1wXUc7RyhhpdQa0nsJqmhqHmDU9vDG9gcWozR8ukzCgtkdB
w4BedN8ge+wn1Sx6LG1fBubKQk8H501u4TsINGTXZpF+3zsxB+SLrDlnsw0YcOvc2tAF/8200hvq
uQQnRiwwWe7RgxOX36+Al9TkSe0Pdt4QIb1Ktk5x3fvga32xI9LT76UZaqGHyj7I6+OHpIBCUzwy
150wcJGi6+BMOc6sQI7/bxiw3wcygKiHtPqZlWatORSGnSXasiFdQWGkV2/JBO+EbNgiXjgtTaAH
uDNxkenWuxEI8EoEAnwMjnbA0NZRuJvN7/2PLvmB/0r8jnHGutK/KzuN1OSRKe5Jcf0a3ZuwgVqf
DMCYEqqEinqCp+id3X082sEgf8+fELBqiCJUm0BTVG4dOnYr0CfwvXP6Dwvo8AJI89pA3aYMt87v
ke5Wj8LkNjyan2Es3fl7C9+XMllorRQfqUxu00LY3JffTM5EYloFugMfGDQoacaqq3XWgQb5xdfT
gxPvPaBshzG+7mP+5SHgVsL5pbcj/JBwa8AwT9WFC+YatjAD2gUygDlUWTF1GA8p2OTt5dswOozk
lkbf0mN0OZ6vnmqIgVi+FEOwked+ke0+Kug+Iw05XZYeO5eAlPfNkDq+MUGQVzIUFtIidcjnniHd
7O1Kx+9DvG7JjVXJzOC7uU//FdXdM6Vs+ceD24CXGOspkAD4OPFiwvOlpKEcxzdAMv0UKBkSuA/e
XVj5IrU4YLKgrm/q7I0lY28MK1FSbqRRXCMpmQCY3S8XRqqJlW7MtN1Bv2X3BLBOQy2s7p9cMRmz
zX7AblVxJWNC8Sw8VI73O8+faZFgvRW/8FAxzuvV/nPKt+tBNT3l00xHcNwWIBFA5ZRiYCw0CwP0
jKCDOodyw6bRWZkYp41LTzjHTdJjj4xCuy6UjTmUbaC1S1ERc3gcz85aESLK85aa4xrXJEoJHmUD
XVxdpJjRci+ZK4gIRJ1cl4kRQJgvhDoDqrvT32qdy6H3RoI6DtlQYlgqKPv+vBwWZ/kRGpq791XR
H426UMqX1oYrsrdkaPYkO/rojQpLvjfD0TLa+y6VEch1XqFXY37eiPFLJWh/a5Ou62JHM/L77uct
+qPrBHgQFbhvFI6/DPXyWSHpOFJZ0ZFePP9UFHpM19Ff56X4/MxrDjF5Oci+9AQotVFxuZBx0Ti+
6nFlj1bSyvJe0idDvh41SVZ7Z1fcYi3hBn4emeHalCRJ5a6kWmAo0EGDuIwuBc6ZVIHQEgdl79M6
ShoxY1UMWPf0HOhsbCQSmGr0LfK25S6App4vLgccqbD3cAZfnAtI0kcYTJN/dY1KNeeBZ9YU8aoj
mELZEHpy4PmRRACKjZvn6IuOlLZoNMncldqHbwe/9gersosunQmJFX3V1hGLeov2IPqItPQa3CkX
/xCgFYIX6qL9bdp9RKHkM+JmUmpF/Tu1ETpv4aqocN0bj+Vi3unVnUr/o+3Q35uvvRqN0s9CMLaY
nv8taGy5f466j0uQ7slGGnhyJFxC17ZjXQgNxrfJJKpcGCR2ZX1YR8+XYzuX/6Der3X76R4o7U+3
g4ZEx/p855VgPDjpkFcRZztIZPJz7oMrLhCIJN9XCYC/lN/zDdCy74n6srYYN7KROnN99WqlWzEQ
8hEwG3Lkd6glpv6di1XuudWOQNRrsj7UA+SQd6ViiHbSDeYXGbbOXaUHh9D2z1KEC3y8By0zGBNx
OVPBYKZsb3/ojKaKkx6qsxrwyaxJdT2CB1bshzH6icV0jGWddyKJr8gFb7H+7qC59wemgf7SXb7I
rYkG4cD9rBy3TQfMAetirCD8f4VIjsGZUHZmKwrebAB1kXw6LGz5Cq2rvR0kL3y9QgKhbrO4U06c
fgI8krP+AZ1xtu07xZg7zqFms48hxYQcDR1Hu9qsUg7Gq7dGBuEXxoz3ZIvkn3oMS2WuNgH/XvIW
VzK+OX9nr4x+NUOiMGupmDhJD+Ry4wR5IFSkm7mI7EXMHPozE83vGfhw3YiB7gYN3kaSwIVVpfqg
yPBeMdeJJIKQcV8huMi1mkfK/cmgUJ5ZUWXR+Nb3PhMRehiDk145jnTLFVI+mGiEtZhOK6mOzy3t
4IsofK9HVfpPsnfdgwD1+Ji+AM26WW/fMEdjvGXzR3toLYSEXKMVJ2uarfEKOWfkRSyKHMG2y64L
agna/SFOjtJ24N4pSyXkLaZGAQkcvmkZqPSaHSGrs8hE0z5UG+6TY026+Sdrkd+m5SLpCa7501gu
b6iO9IBo7WwgWsC85OQ1Z5q8Bia5Pv1ccp4RGn5k/gbr8XG1sVi6fneoSjscMWjcsLayDI6UvZBu
FFI98xLOOSuZxotIKtOVqyi7T6xpPt7pUtJdPaqwWPQiIw3RAn3bOI14Wojn3rgPn4uSJr/Lo5QR
FBv6VXhC72ENoh2JGEsyb6lSwyL+g+ESvqGAG3/xyoq0lNMx7gqFJCq74TtBJTeTZdhUQLSoz1hC
RQ8FAOqxe+l+xIWUjGFjOEes8cBzNoALX5rBXB/Jjz5d2pUvRInAytmReKwLGoLQmGbbMQjsMhQW
g9OWMhqqfQ5r2c6qzmTeuwZju23OwPYvnCWO6RxZ4zfW4vupWy+TiAGYz07AgXZ+k3E3pgC2VfPZ
pl+PlTupiR6505m4bc2nIyDC45Pr99M2HdcOt9Li9gk+bLjmH3qyQaZ4mITzZsaKCt5PM7gdKm7h
QoHNfG1jzLroj6HNlnM+fshXKnqVIrY1UxLoxjjuSCp5D1K427KbIuBG6lpLJgC2DFRI8tqIwSdM
u9GW20NuVR2E9Z3iVZZ1oxnJldhXzNF4zoJo2RtiH/AhUFh2FgdGFsSrCxw21BPGwO6bcIzzdijv
MTuNESrXNGMaJZcbMeQBfhTRELl8yR/mTbnCiRwnTjrSZxEYroHb+1Z5SuGjX1CiGnjKXs08FNUU
4bf+8ZfCdY/8YyWTCptzA1y2Pg+1SJHtWE7JooC8FtSWATyY8lFtdxTZSfufA+kNpAjR5or5MUYn
G/QUEoz0qeyDzt7lG3PDJGtVHlLS8NT7nxPdv5l+kfejpttqRSmgWVmbhgHWXbddh1VuIkPGOP7C
qIUPLp+YKB2h3wSrWfKLWlmbK5NrPdfkhZd/XmSx/g2KzpokFMmCT/rJMjgay0knie3IK4FyB7Y5
yEal/6DYACeRI6QidLIgnA/2qjdm16cabHCzHy9RyrezqM8vovuLMnHWTFMpxTCQlMPzuFdiGwks
wrzOjk8FlnUupriOzSUt3DpOvryqh4q1PGQ1b9NZ3n7YqwJBtxzsGn0rzOP9ojJ6VPA+dVzPKGIK
gIniD11SJK/poNgH7jyfzkhdZye5h/NfzAhBp3gTRbozFYsYiA2gXvBFZ2i5AxSwaCEcfrZ/WPWy
NT8ddbeYeYacPpuHrC5yWCJGB+p1rX6fwhDXgpf9DNQgMIlPiNAOjSOPwwMLC0VBalDx0ESEe+uF
e/1Barki7JGlRpWiLbwhs9aSdoNOBAd7M91hayKqRgFqNHETp34eko3D5PEnIsYOOwQgEFrytibE
0+tevfGHstg2F/HBIqM6LjA0+lfuUOd7kzg4zk3MR1BpEtUqFAc7PH639C+w796cnVBHzSJGHncU
Jt8/tCRzJogs/d9OAkLrIShgKimIH7YKkA6ayQZ8mncU5VGQ0bHrgUklXCn4kqrcy2LfrCLWsioH
4bv7n+3f5JbIFX0H+UrLhLZQMJ4KNF9rnfHiqjmTWtxPXYz0ROhYcBh6M4XYppDgkCt0wBsLNb5D
pNoCisNFgQy3+NAGj+MUyRXJ1FVdTNxiyKuovYuCJj7tN8iKb912KtjpwIONyOA+CQFOEfmYH3jS
eJB2br3i6ndJ7Tbtfm2kz51xVz0Y+hJLuBzYRiAxzO3HWGnewG2ZPU+mvWycpT2GPfqdeU3UNmIz
QQIwdYbiTk27Ncbc51OvkWVFfPju6OZ3XtwJFuD5LY+G2pjdYyMBLxaq+m8X9AIUZYgkBSIKtV4o
W5O4JQAJMlRbgALq9d1v+5WlNVGuynInm4X2wGFTdDWEiNE8WvLkqddIb8e+03orE4C3lsftde2n
KPtEEa/IEOtS3KdVmCcDokFk/L6EZym+b0v7kf946pghORzrObJotIRYQPXAaB322IiajWT6lBfy
N7BUOjFDAqdGVroafpA8VPPDmmOleElG6WvU3DB6f3ZEt+NzuYFqPSEc79/d5o8/2SZ8IYa50JP9
48V4UzgczmnSLv14WqcoKHJ4HomrHIKWnVtVBAyEl2OTRppPoG7/4CqqS6G+pZneGsuRS8V/qzT1
QBwdGrpso8LP6iFoY/bVGpIi45+UaXjmfmPrhS3qBmIpjYBBlO1NbE+dzZ8EUa9nKWcsPGap5hWO
/xLcyOpWahEWo+sYEOMv5j5kRt/O+6MnBcKVoBZ+8XohJiGcQzfdQ6gEK4mjs6GSdpvh02O6q/co
qqSJSc2+/tNEBjA0m9I25xHMcZKlwaGVhqK89G5BzXQvRPEHHe2/bW6zKqx55c/e19LVGCfbGskP
isK+8wE97SJXCOuHkRmnLm8f0d3jXO3zMDi1RD7a+BzFLRhY/pEkQK8Z+u4AvtYh44XI4FXqRDe9
cXZyVPif98JUhG9H/otbcgLliFsgc14ba709yDVFBu1jiB3SC/wbdeRUvAjCc5tt4R1SoQn6FvoV
CRDV9ZwX0HEaODSplYx42AeOhVr3/UsWrs86hV+T4egN8qYa+AFLRFTo4fISo0IaVe4RZVd+N1fm
PXkWuV4yG8xrldVnx8z25yAh0s2xJh9ImunYQc3KdU1xFdObMZgXxLd1zXpCz7WLpO9OcBaBZQZs
8mPH0JhJNDIdhGj+gucp9KiJweBbZukDwS30TofIiT2ly7EXQjUWhQfMhrmTjFLqAbpojZ/6/T7G
pyA2rzO0J9FlxtqxYx1I2pMofrabq33Mp6ZYpqQSrN1y05UFBOhEvf7eeMZMZ1WVw+RCV+7DXaI9
oVkrFvM2+Bv7r84aU2f2xM0f95R+rTLgYxYbfI1lUsNQ4lexlveyzhW2eynVtAtnIDZa4BhwLI5c
yCnyh8sw61hE/x6n/5fh9Qvbi/IyHJbwvZXf15rEmu2nFz3ojMPfwGXccj30l3TzbbnE8/abg6VL
prMe28lf2K+2Nwt6OXaxTEM5ppULM7KTJNnFXwaSBG9Xs1R49lG0qe6NUPerpnstVMno2iMCpyT4
FcmYp6TWxtFoJmX8tU10XqxzoYlBXg5V8q9PPfEw4CNsAq1ROdDLFkaJyP3MJP5ornv85u3jXMiR
RWVIf/dkTa2ks2FsbGvlHzzchNqNGO9D/GMhWbs/Hmg7CskzkYDnKVZJkHFkifvtCzfLVpCq2bjR
JnbxTo/3tmwgoK5N2usSUnQTLfCyngm4WM8M58txxkh1X3vh6GMvNukv3UtgoCs1wRRfqSNAVpvo
oDDt61iH5acw/S2u0Q2kfvkPtBB3bgfHw/9xDRmqEJezf8jxsL5oii6eOb8bcjjWZnqPSRT5GPIX
Yg2AHdgQZzBcvIq9wOxfO9sifyK04/KURwC24UZoG9erUoBLL7Ca0D9DOck6gRhWY6RFtUHOpdR6
Q0FVtM46+T6QTSuDlccCfq5k/D+XAlp4qFXlG4TfE6GRC/9kuZXcjt3ZPmU+X7eYlvplDbCz7gwu
Wl2ewx8W3yLYpO2rQeAp0q/uuifJxUXVUchqhDRz/iCZM+NdjIjWH46F41Xi6dGSchP7EfwhzVmb
YYLP+F0CgR8Rvh7vZvkg4nc+/5zDEUNkxqiKVjhGA5ANnraxXzXfk3DwKAmyNt4s8LPcyrJeuRBK
/GoUAxUfZh0Dwv1/wOEC2XQ+SlEzGIyMjqI8Roo5XkI2VhINXdLt87wKnWTzvFgoIz4Hw5BZjT0J
r5OhWqCAXjSiTLhHyPZwY7rf0WHzVNgU+wHzrBzy/3uLCFKs4o7gacRLtWeFhK1as4VKYhUjP8GR
aX4BJKmNPbvy0P/1bfO+31l57W61WPkWffAQ0U8zjnhcEAJP+2K7tBJyPSw0TwO4hbiRuU/QkDUu
6iQblqUl+xuJAGxj5koxciv+zISxzcmKQPtrjHLJCC2aY83DN1MV4r8qcPrSuhc7pbJ4T8i+nQsc
BgfWnd00ZNlzsQ566Pw1BkPY3iwvU3kVs4cJnMxMvoJHBcrQ4oMVFvlTAQorCT6XSw/xxPAAMCb/
IOira1k4ljBm67eaYRRClpqjLQ1FQ+BylXQNzqJ3FbV5RjR/nLLZDVtngtPhLwiKOh8H2PHUpIWB
NbxwIWckZC3jxGwekiEOwaMyX7iFTn0BwvPlel9j25grVLRVB3vhC7m3e9Lkl46A4Mf6jpOcyebC
d9QoqnqrdYO475nA/sC2HpOkZkkv2YvxOhHSbxqS+ubQ5nDswG7cyTwERauSHRd85E8viSk1fL8e
jK+BlJm/Fh9fINtEFKJ6IutstwmSh/gHuwMm4BBLo609UU+Dk5wlhQp49gRm8AST10gm7QjR4RU9
eTmzX3LRefOchRzu/9g4VplDZHLRbW9y3UdKdAEgUUyqyCoot2F5nNoE0DGLPm1ZlwF4d5WI+L3+
ctTUT6SOaGd2QBhMB1iDvXK6usL1NwTTtEukP/S74KXS//edrhv4yGXQrU4IwErQtGT2Su17e9dD
qqxJaS/MrtZB6pItokw3AQcGzMG7gf+Yq6jMPkPJyxqfDmL/4EaRf3U0c9voV8tNvCt6+aQZhkIW
EVa06jMwdxNamRluc78Qywau1BEG4fdF5QAUgRNeq392956C5N3sR5D84037QfDBr62j/Or69U4F
6kSKysgfJLbVrrApNlT5AUKohqJG19QG7waHErn98p0oCq63PtN74hQWIHY7Gk3CHGeut3mjGZE+
QeQq6/jUxvyEFrAa/cR9rGTDSeNaGhZGlvDNS2kPiY7fA8HwuHT7uk0pn0rHFTwlgXY71eO/ieUL
aBs/1EWviNKneRMnpIPWvGbESEdbrLn0zEa0BjX96waKnfjMcYZEv+JkoQXnMn6zjaldhiX6yF1i
kqLKLr9yUPYNQR6MylW+2DuekRGVTx2uOflcIlFXtxXHxc+bEBKcDKeOUy83jLYat5rl9ooewvdQ
4lewX8cigvP2G9Uq0nnoFePTcelZc84GH3/P8/PU9oh1F9+TbX0MsbAzeXAFEqNCwyqWBbiwzMQn
GYGm39qSRw1tMWa7OIyusOI2rtrDX7z76fS9XPbiDdKdO4Oty/YQK+cQY3tkE+y1Xql6EKDmI360
OZ5gLA2E9Itdz9Aqi2oGQtFDAne7TqfaWRxKs1whWclh+Lg+jAxvqYG9CPdeuOSOUkCIG6doTaQN
yEIjrkOSJ1WUhwpWYSqoYMKw4h6zp6xzSwni7UIKz+hebm3mr9QKZDuEN16V9c66lQBuwsUUonrb
MVODv4TBjzUBzy6y4ubfNElsj6yeDPkXGtRWWpn/udvEW4UR23eG1/JSlAGe434KfD1Qe2vFO1JI
1f1JIueaL0H1bkmIdzPM70LpzDJ069Dp3fFgGpWMY0mevi9Cw//nl1tdzHJ2FaneKCKcEx/++RFK
oS7At4zK5gdgMQTFVeFHkz+JFyU0LVkEARl0d8MykZhmWgYTkSQzSIPXavfJ3//+gCDsAOFLeHd6
V8+KMvNqSIKoWkXBwctfLbf+Wu8nfSAK6ioQe0lxWq6AZoAVp55Avxfl4AwJFVSU7NtJqYEJLLHR
YPzKMY1sNSllOEPzYe6digw9rQPw+MuJ8oOvq7LO2cJpCEC1Y7eT/BSRdV0J+mZ+SphBtRRDFWb3
f1FF7Z9ibLALns8hRLSoU6+HFTN3vGkaJDnNfrE3dvBCH8hrGcFMHOJl6h6sWImeQyuAeWwdTubC
C86Gn0bqUQeHZdc0MBPxElvVxsDrySFojJfr05itjS9dNth/+eokBHQpVJYGckLWx8IR7K+Tpdve
9/SWdRY90CXP3bLdPIN4Fvksr9sMqoqbJpdHeYKWb17wl4L171PtDMRR/E9bImv/ofL8l7DhPpVi
NSAavlH5gzJGJoQlL3TeeQIPAK81KzVTgioDI9UGHUTY0ON2vEz0LlHytNU6G3Y50zErWR+ubuFX
C0OfOMNa5OWVdKjsCvhjSpgRFtIF3GYetE/KvhsRSmcPByPJ5qzXzvLurd+JLsOUn8/fztlc8EFE
ssRYnItjPBS/HEUr/Cm2NKkKetNOrWjfBAwEqhWonrk8/zGVo3Lhs7m7XtALB0ZJCvQaF0BWFUIj
PtF7JJFy7GbiIdhbeKKO48jXUdEbcU5tN9wMjrFKj347OHD3sx5LEy80BEPMzCCO10td1/Nq6I1r
LwnO/yqEoTrPooySrTNIaVzacIe/h1KOzsX4mH/IAn3K0lpcoJ579boBfEyASJ1JkLRxz708EJnN
fNX5JTiF4DoXIgJ0cjUxxejYVg7C5rD00KHPPQ8eU4u7O3G3VUphofWxGbTJSSRg04bM2CCjjNwV
8VkJFgPEowSJVTf7iCKz0SbGlu8zxjNSlKOudIz244QH86EfdIda9EFXYs3+WIszsb99lnzqIFoW
NH1AUhb9d6rTAQHsZ8Pu7goReQHfs+5J/5sxsLPgQ+ZJP/g4aAgiMmQipwH95vUVRuOnKzICqCPf
RR8d7qYQ3n1llsNxcd2JkE3FACBci1pp8dFDzZaqpCk3GkIkkDNWgsGclQtMtRssdpHGVQDZ8IyN
LhCYtmn/VlM0BJbSpMRoKldD2PL6fJM7y2HbjhmWoDVuqEbFXQ+B9LmgaM9s3CeByFMqSensRQRZ
6Je/Awe7gxnjQudT/4c4z62HOIGVPt7HZDc0qFJX/xYh/nBfvXEZH4lLrAGswVUv955Wax9vD3wQ
l7eTFhGIkpD4W8iePqCmp8FekSJ+u1eKpPPJO+zT2b3XkitPaorNJ52SfQxnNdVAK9S1N7k+QbdP
uM1OMeFjnU9ETxgevf3dDd3MTRf+owH+OT6O0Izc4d7/OlVWdXZC2m6aoJsLLwKYCInS7apJtHXx
e+ym56W8QNyWj/B6VUyGtb+MmLwtBbeCopbUXWagbU9yUgZnmOp2XO6W6FhZkTASDj4+/RIgZ6li
n+2+bEJBJiY8ngzbisG+PGL4cZvbdsNWIN8EwMeTPb2M8tI0UfWmb1rM3K1tGd8zCz03H49OjFPe
onhaOb4Logcx8nY6Z+0KikEUapaWOrk32EYI22uE181Be4itVqZOCnkC/FLLxapbzhxSlsdkjvn3
xjzfCb2Lq4pU1tRj6+2Q0kzBYLv4+g+14UJ4PJM1jfV/aNk9j5OILUD8wImCOVb4Fd6kN2vQRadx
wWmy6ydQQ5AcKPlklSRqVYqbEVsXTb5R46JVlfL8OxKJZh20zwLOMPFsbxUgnh/5exrKosuCiadN
gjziHlPnL/4HDPJc8drtaiccZRhqg/fDJ263OD8HfgZ73lqyxZq5zlxyTB2Ax7q3feR+hubRmynp
4MLfyCaJ/bc4YsWf5WtY6tkMLNpyFnlKJz7sNzknc+WmGTc2Xrd56eSdayWiRQTGxxHLdwRw6jTj
+O18qee6i1u0baCovZ6CfuR2nktZdXhE5/CZJmpMUYBYvaL6wCn96aTX5EjgJPDC/eCpAZU6QuGB
f9keoG4djjLhkKudkfhqBRRAlLiTyLEZ3BtYV/YYvIe++IEwXsstbhSrumWElQQnlqXGl4hwQ/YC
aIgTQCsCFPtdCBYpU92HFKRvmYHsP+xmA8EFz7xwmaqgZaklSPwvRHlesMRU76LHz8BOiyisImov
+yGqP8FhA/Nw8DprVA6zRDadVYPwhLIaLdnRsjgd6/WEsUauRAkdK8Ctgp3eZlPxhfx3HwJspiaK
fh0d1twA4Z4hi3ewarU+kuY551+em1D3cpubJQowBp/VE/H8tAJnEMqFNbVCALngzP891NcoX1bo
fZBYHfGomS5Y/vLL2LEbImT5GwP6YWISBsrLdDunfZBFa8+oYnwPtce3pZk+AmjKKffuIDPhkRO3
QiU8LjixEEbSCepo9mSWSEnMQC5PQmnXK6D4HAJ1d8+0vJyqf5EewObVcgrhH8dqCLg30l+Y8UUO
lW6hSDUYRVUB/B8XOS2vEcF/cv++qmjphMRagHSGQ1ozyQ71ViJQVQtb+s2IucE2Rm8s4sXg/ASu
LmhGTM01OSfIRwbsjwTIl9AgHky4XfOIeeh6G//gy2KGm8LpdmelUPCZ6gF1DM4Sa/SJbTMCCRut
Di4ek/0wQQayj++4nIUKbKGPaYYMi/uG/SQl48J0b0uctCEKpwVeO6yJ6ZMCrvWzzPVfPNDAEoIs
8OxHcyW3S3mm8iK1Gz0J7oqb/Ch5DuSikQ3HI5pDmvlleWl0jGmMKcerB8935xrkckUnBF8z9Dhf
2g/2mealEFXnHfJO11dNpemJ6Lc1Q2ch73bupqnW4fSuyCoFCVHeP/nAHlij7VQI8ZWpHTHU6y8i
LI09zFoeO7cPTdyDlsM7QA9t9F5m8TVEgXyrUiqrBLx/XBMz0Qbe9Rv8A6QQg7xNZ4CO5Rw3ZXOu
QeECSvRjgxSojmy7dc4KQylm5zLALOTH4qQhTebdRLJQRsFzctq6ZKkUUpuUvknYQHk5IqdmMhLa
d4XJojpIO3t4oRmbjlJUAj7O4vcwmoL4PMlwE9bPa8ogrQmfP9IRmaHEqqwD9yDXwVGRntN7PwvE
hIqE4FnLh58IShYt1BawjaKgvfD6+/osuw2g3OeWvlmm4BCLKQyw8VWQA1E1FQGXbrPtu7eBD2QM
HG+SN1LrR2su+hVIQ0IHiTj+4iQF4TTEF3BLw3Em9MlSZQ8MFdgaQ4W6V91DgRt2LV1kcUd9GWvR
ceyDX7PWRRapJ5Gu8jq81tRoKAEt1iwKaLe4zSIgdMkAUY2HppXwHBSUFqsLP7sXVUrvQTr7Ldgy
2ue5gFbRhCjOn//J7RSaWGrDnXHM0ayWNnZYvDDv593c8v2zNeR7MEjnBehRiu+wJP9t9ZMTEdRq
7q5OpXNmvXHn0I4CA0tVU2srOmV4slKvAe1Bz2jfyW1KjwcrYqEnW4xjHK9P2P0fATMKgXM1T1hu
kVA870LRlgbd0o7zp3moBbmtNR+iGrLjbBFtJKrFXflkBLXSnTJebQmJFs7osDsruyW5g1C9A4Ku
IB2hOj4JCoic/wXPUsC2W2k/uf6OcD539UX1U0MtBfRIHEZ7ThG+VXRJ5mdA35vKrzi2TmWVswFw
p/jRQVONA13Z15CAkoXPTrg5zNE33NusqrZcH1gSx3s67oL9hfoKf+LcPZiVn1RzRHtgpj5EAJ84
jr/GwUySNBOu7j/hF038LfoAqbR02iAcCabP72Nz21F8umdMsLPLADFNPK9JU6CN4p46YbtxNpKI
u3r6EVKVstHvJjN52DXbv+/9ygaodJVrz6dUc3QlLskqNx0CRTRzSQ++VRizxfJ/s1rdeH76Z580
mvUK7LhYRuCFDlkzGODZ6OLZJzDeY7jS3uoanGwU4Gp4bah+P9oCmgicimEzIJLYcRZRDxk6rATS
e0D79U5qbNg1NSpcpiz9vmENszgjq6J9M/TkOAf+6YB3BdRNmxtdZC2yinHJPZ/GKI/kCaoaFfVE
CdPC57yNsv4wtj7pwra9mTaqKYk5+uTr5ZP7gCQjRpug2bJBVvgq2QyXUQgWdxKcdlH8VwV/d+L1
EhfZoG8MBiCc7rN4GkDlm7rIoKYqAUqkjeuH4LqiMammEaWiZhHFIe8a3RIk0GzwZfmvIxRs+/lv
w2Spjb6D1U53iJAwHdwgnqt6T8TUN08qPqn+KJoHXYibUAf/EoKhqEMO8VnUEf5UJ2uUZ0o/Xivr
hRKnaKbJ6Nn3BP/kVuzcvExL2mWKVn4r1XpFdg1jnoieXHHuic09GiBNsmevjNLWsMH+sQNQ5fY5
SiYGoSTgoHtfbIbiW5zv0QLaIrao6loo3j7xzZ41Kj4ffAo4A9hfT04T34xLSRcYOtmgCvfpNmNp
oq3STcc9FWNV9dm0KO2Pq3SyAO518YQ65tBoksGedhtA3csDoGXL+HBL81Dj0X9XAQuAwfzEr54i
gXYHQiIuEjQ16xL9+fJw0RTSPOeboeYgjOJ8cZJauyjOR/U2u7c7BhVfaIVbTOuzdCLoKkt/GhJX
7RUzOc5xWTwOBMCzDTga6ARbA2Pf7cWayUbBlduvgIyGgwOJPoyrIug7vaFtWcmqF8Yd21oa02hc
LxjPzMgP32g99NToEODzn+MGQcsDfJV8SIWfsGHHwV1Qaf/C7eIeMtHTVUdjR6flWUImYZsX6x1t
e1D8gZ8qKkFoAd/6QJ9NN9RoHgXDjIhK08M862gz7ioLPyAQeHYffdjXCW7jBr0qzkzGUOOFyHEm
/8iIuFxIVHdAsTweuFanpSXmFVIkU4/YiJLbCMALxDJBwEbGYiYLaUno3IaedGSGH4HgwTo2Pej2
908cmJYO+aArj1fGw3d2MDznnIGicSBJVWQlCkr49JozhBB+PPvLdCwQw0AZxcFhEynaPU9+y5Q8
4ug+zzz8A7v9vMnq02W3ttPi+id5+LoTvK864SzkniMCpcAJ01LnMrtwYZdRu0On0XOuk/O8kvBx
565qM6K6yU/xL9rbj5qPB5KONu94dyt5KNk6z6kWXM5IhVSbWJUJ+l+AcUqWOLqNo+iMee2aC3Vn
C09JxuJB8b2K2fMFKnbqID0Kx8/MBLc+BWyIQ0k9infl+1ldSbEwwQS+9LPkGBnLixfz2P5anhoo
TzRW94NymW9eRfM/GhzF5CLn4M2Ke4Up3oPblxc7lWk7aYIpeCl0JOAp+85QJczlaAukKUo2iYbP
7OmuU8s7zrsyV5WMvhiIYzXbMUQp1xxhYfpLe6WSunJtafZLOBlF0i6qBq8ewj+v8pCI9j9Z1fNP
4bmveQ0QpS+I5abPC67jRMQf3VDkmv65zjMFjsSYxVmshb1yRrMUT7axSuntq8sse8zLXE0wCX7K
DqoCc4vAA0CuKTjycgEDUDuK/cQMowVSiHQJYfVc24omoSP4lMZyxjZN9DW1TU/2EvwHHOGHtFHJ
y/cvNFPc+WU8d/Uc/tNKvc1VysJUZcFvB7JxEF9+7NSc2NUf90M8gf3RPjgVcm5rsO2JMrZg/ual
PnXRz4kp/sOPni0bQph5QKauMdbng4FV/7KzqrJECAzGekXFj8Cqvb0XFwqjaFdcIQyKZbjSYebA
TqsrSjBvhpYOBEXbyZxGRAQqd/SHxPrPDhStHry/wPVFbIyqpppnTq3O+V3qSSgPmx9XnaQBTGIU
ebAbLGAv1T8vDo7RXY/65Q8SYtMDK992cadRYL2NEXA7LFEYVuHh5i33DMohe+YtgPRAOXAAwW1w
7v/4vYXNNYEauSxbzLQEGnZYkYrhczFDiavmLjIwC6uZXTB8UviSIWbFndSsT7rMEFezTGqfrdhw
XyJmJAq/z0VSZkAW4r8S5EtRcbBGq5LpEZVlu7yEgypXTx/CFYFw/qSy/oanZf6G9jIG7xe/3Quu
N+upIvc6dVoH65CCy8vTgJA1pYlF6UUiOBk4tACOM7lEMgVz+RVkg1qB2rz3Cku4CvEzRBU/xYWH
IAkHuHQQFJjuEnFu/1x9bepJAW7bhSsSY9tO/mgUIN0YhEmNu6dChb1ofK/r5oaJAl0UReuxiRiJ
pXWwrH0MlhEQxLUggI3W/5mX4OoimWVlH7v7fzUE4JaHZiswz31Eumz9NQVV87MI6Eg8uAxvuMHb
l3Wcvh90G/WGBJIquwkvo/Z2CFAHPnT3E5Jx4whip53b1RREzEKBalcDptIlOsSF4RScvXv9J9bx
4CJXxZk4Ci6/dxlwg8XTLA1aIw+JQvMX6ou38EVkXAIpNCaGidOwjgt+KQyGHn9jR4hUPehJPziL
qzcCc+coSK+690X2uW9RUI0dGQsWdArxoOipCKUPhUxenzt8GK6J4d/TLAqbCRXSpE6D03CG8OxC
AmgyLzfnDyQ8ukqlJVkExZ6LBY4cC6uwwzdoOh3lwxfNMPxPyihpd3KBdWBZpJPn5htKzMhHl5Jw
z1UHtp8HVVTumPAjK6pGhhuVqrbi9uAdItmAVUrDzgnyYLz2ff361dQGTWEZ+RdMHLRAubPxrgli
hxLH1r/tBuAePUuXAEuVUT6eWx8sYTJDz2Y5fZrW2S4MqH7lvUZxGSldFbpj9+oMX62BC1s00NsS
7UGvFh7dfBtyGTqpUkNnEHKC5hBjYsiT/Ax8kF+SMr7SVgDvZ3627xOAxyXzI5brKyrDzmhua2Yi
9BVOqj4LFpIpVbNSUiErKzip6CwfYSF2vylNXD6wn/PTreKsY7GAdd7G7BTbs5Q4DkGTDLu0554V
F5UQsMsCt+Nxk9MrJphIwTkbWyEtMEggXfGl+godZFcByulViZ+Og35VroMffBGW8CRggaGR2eXc
gnAYT1sSO73nALwG+ZLJI0gA3J3hIHkx1wSOf/z3/utzH/IBphWU0gfGX4IaQwIBlXfYu0eaOjQe
ozot3QI8pEwAkldQDbVVgi+g89YzydoXRlqeVDOtTsitiRJKOlxVrSzAsVOsNWWmYhr/Tj8w0H2/
jPRarMTfGHk3t1oEj//csf22ab0J1chIPGMhY78J1GQyKDutAX8yBPIW5d7XhfSeB7pmsZXCyRyb
jSMvfcgVgQ6KCrNTglIFfysUdcrHcBWZ39xW5toSaabibYntM9XEyc/xP4OWvZ8Ko+Y4fdre4KQr
vDZczsr2yCRJTUoyeAOGHARQQ78tk3eoapDESU+kI4yFRoFcUqA0AdlmICTI/S0UZqiMIsRDddFW
5oDMc9PZmGg0act8NpLvIKjVMjO3JjCoz2gnFUjQda7huRI7yvAXnkQRnpN0BXzy0ukO9CGoQM1A
D3Kj66wsRr7WMlnJhydOAWspG5v+4ybfTcAlLOBR/6DlBrBgXmDlYda6cTS77wTYeOX2svMqe8vd
dJevJES9mp8ZCkQJvKgqrnKtGNCaudsDefUFznsCWWHeVgIQNdgMOeVWk9uV8P0Qovvu6tdii/Fk
515M0omdERHvSf/3P5KbimlsZh0gP2/LMOhM+YHZZ4ikGCGouOSNZPVFqAs6QcY21APnkOxEulql
mbnAEvkwNSEwDr+R4o3XdsvDXKHCxPv48lf4bbHmuHsX6nKeJTOiEXljedgrisGNq1IVEJGtbPTZ
ssQ/bHWsGibxSgg1t0X4KuPW5ByOro9U06Wi98fITubQo+u4ZZilxV4klC8FNjdEDFq1x/M4hrka
OhNq+bfBWC6jk4SPHm7ONKU76XkaoUx0i1uS6UfViudPV+MKyW4r43ic59Yh5V9nThSoluVAxumC
cGWReekLjd7z/N/Pes+Nv41nB85CBdbzNwy15IDUTpKeB9xszIFj2VvBC6AvKwWEhGJoeQWZeOoI
OIOwdSK+xclJnSiktZ5+42FMkJ3O52pw2XB4e0M7U+aUAi2NYU9PFiaExriobIfkNQuMvSZYcoOp
2JUHNHASqs/MyiIOFBza6NXPEk+jhrsygRq+7+w3VyVUUx0kTzZ9LfMekDzG1lNntyGVwarnrACv
zU+J8BUZ9bhLxLnemJOc5rxNdOGXJXHEFWv3VjZThBKEllDj8BoGmyVpkvxUEwkkf7/DE5GpKlzI
G3/kXjI54NCYvzEnuIaThY1eOoU6uRYMtGqmOWDQDG19Z3N3yTcOLl3usjkdNrEREI6Ps9G/LQRw
RZozNJU7qvbWu8pk47+B0PXWq0qncYUBdOK/UoYPuZk1xiLc6+3nvslq705OI56ws8QYIZUwymvS
WWs2te6+T/eHGd1HccEtbW8tMWuKO7H8ZVjLh4s4atBdd6HvyD6FwycPKuqp2hSMEhmTmmIijACZ
OyfKDV1fdmPn6jYfRXPzgrgy/cJU1mc8T2LoNGe8pt8gE7FZPwFFyd/lQDzEyN4lPv5uNeMdVYlP
lQ/QGKb1OTXirgsPr1Cn+iIHu7dqLw2hvRNigMQhduRBj7tc7wZsDC1dyWE1+0yd31e+Zs6Gqnwj
+sahEe6hi9tG0D5kXFNvshs9CK7J2XXGWg6EJ7r0L0EHcvSw9v9ZIZecTtD/BNVFTe3vY6s07YP1
/uaBfqE2eDNuuSSi/H8+64XOB/EpY/vrvGhmGizfCE/b2ZmBDevhw+YjEBiPwzeYD+kNZk8kyEAP
LrVL1ypm+NDwy+ElH5tiY5fBUigw3h+YU+RwtQKUJ16p648HJOPmsrk3vafaZ0+C6FpebwDL8ZoX
M3s3K131gOe0aoAAljmo5qwuIrN4hni9NUashpASuP9rx/21YGX2d4qlQrTVk0kxD39NflNkETs8
3qKj6YDl32O+aEoeroi2KX8TujzdO0jhSOoX7jvOp7/43HmOt7bAAPIDBxExfyKTrXWuG9M/RPnQ
NYGHgSc+poY6ol20zayHPJNGSFV6rfwwR4RNG7OreZnwpI1DliI8GZDH4ns1Bs8C6IGV5pfhNX5b
QdaMVpZBXWHXOoDtZo7JjXfZgOJqPHSUkKDDKWyPbGWUWb4TfQdgmIgAADbJzIyUA7nr49Obm5Wy
f3D1lpaPJjseT2Z0ax0RSl7pHJhSJDV8i58UdskwrwPxFHaJRDRKg8NfpCBYtyz71+SmBBYvQKaI
CC2ZxAI70Oe/7Z0Mq4sxI/uy0jJXhcVKoyVUcJUKmepP47US7mxhf2NOuyP/M9Wm8gASPLV5t9pE
NToCSYJVjyan8zoqMz16JuEoELr8xyw7i/uJ4CjptHZIZw/pR+UU4gc+utoaxDBrYcoYLelOvdWF
3dMxb8aYumPtTa4+6UN5tkJNkGNW9+YUEcdiywp9nIl0XM2qtLPYDXh5JumOJuTJO5am0n4NcJ7F
o9SchyTvRGFgDrgUeR8svTHrO/fFFhyAcUdFn6MGuMLKaZPd2tNHvNlo/+dKDN0ADT8oc68sDY0C
u1E2caY0Wx5YzpDH7WIxFhDKCjfpqSWyjBz9FSzL/2A9WdC8qW6YvzseJlz+YLOKF746vINMVJTq
hBcOUUeThRlGoTUrNzbvas3LHdz0IJuy7pFhp+eyOqe9pHiH1xkJ5MtgdKzpHS1LBB09fkEA1xp+
E+ah0LuPx7obcg6zIDmTrbj6+tQ24VeLWUUpdDrOSyLfUCRDW3Ybbv/9xwChLBQ8MUkJ7m/5N+e4
NOH2dtoVVlxfH99YN6VP+UyNHmFmrebhJG4yPTq7g1DISzmi0q3Hp1G4h9BECcTvNd/nkg+XKVZC
lGrGUR0SLIUAuymou4xzVBTEAEk8Xd5yfzN6VdKZIV6zy4xDkvNE8b9asy/fZcwepKD+bEOKW7mR
/FGRZ+UblmfLuU4zx+vMaN6qdWfX/SI70B+zuAY5N700IaFHUK2Rbwk9L3lnwi45Ove/IK6u5sAD
LHvMVeFGgBmmilcnKMeJgDdn8DQjeQ8GOYID4+Fhqx6HJdahDKNRptsBzUQEvI5h5iqb5pG31YYC
G4gqs5/bljgse3Fm52zV5je8+pGEXZfK5VA564KMyN3CRpenYtmtlGrjg5wy5ok2NX9X1s2wnY+b
iDLGV66qfXXcn2hRUYuyQSeru2vW2/JOFk3DqX4tWCW7H6PFrJ2btTXNa1VKspBMCWg9aMDuYaLo
TxOPnYYCTgUj8wWvIszjw/55PuE/LCwSlREGePJmAv54/ArqRigO/Bc1djQ8+0AYHK/hVI0h3u4X
QtvT8sW8cSeeqSllOcy3CN58QeNUhomvJdJzL+N4DnbvI+986IW8P3ON999xHm0I/IfUciSPV9Tm
DVfjO9Hs/qx0TbrPim/2Xd32uX+EqKfaf2YMk3u8iu7FD3Rk4BJrAJi0o9iCkngNXuXOj2W1jqHr
PrHOCq4qhOww4L7G6IdOtOoFsanhlexfE5D7qf/mgpBQm9XI0Qj244+vMjgJcA8cGxUlRx8XKfi5
ytid1fsCEQmd8KkUZmPcop1PqqT4HdL6FQrOwL7VwVjSnvKql8b9MNtTNW2KAxHqvD7vqGCkbrvA
66SNdbo+qZIEmhNOwqA0Di1PwWquUBko8FjY+HGGJNKB9PgRvt6Co2MfKhdk3jVoPQ99O98qQXi+
MOOlGhjOGHGynyxo8mRu+ztReWwOS0iauSixmQoAfC4D6+Iit2Odwf3SfDRCMaaZSzdR8csaBKNk
Gry5wCgb1SHjXJWNkKLTGqQSHH8UX2/4oi/bAZJszXcUxYv8BCWHEgxBmiq4EQqyb7U1npa4Dh+T
LKMiVdowrH4maYxCDCGTfU7YC48u4OQiZ4S/SYHvII74woNLqT18UOb5OM26dGQk7+7uMM+xAkiD
RQ4vrf6jPiPxDqZjAwCF1wby3OFNust3pYWgdbK06KMFePMzL6VpGTbdBbeA9yxg0BYhxX4FnCAc
dXSzSyMl/4C/tzWIo5TCm/Vq8Qoe3mTJGIPKgSf3dBkRjrKZOBMohBWuIw3qMkYobJ58j+bi4hZX
P/8xMGx8IX+V4Ac2pTjb600eQfizPXQSEBvd2rLR7TZCmV3YMk51YUwmCo+Do1zn131JKS3pb3jx
IXvRBflUjLey6Z4HKjrw5RAnAvJyKwQVM2Yo921RFCtT7oUb7oMzpqwmXsZN3shi3VTFkHMAf5za
+iN6m6smRN2TBV0YZVPkT/aKFWpXaT/kYQxCaqogwcNqD15cCYgtn7uZUGWlXKlIXz9zXT02rDiq
CfH/GBI6O9yYjrIR1czuDLAHZb6u4DvZ6ySCnsweIjVNy23UPi3ZDaXRyuDs2vf5Q0C7Icr06SFi
J/HeUbOv7R+1OFiKpTnWzSh1JD0Xgm18HKLiKH4na1SsJxfGyjotlW+iUVe8XMq57RF/1c1fOimF
CQWY+sQU4en9QGs4fMTRwXWHRoRTmWLKWJikwbhnIg7Ri8l15QZoteRHEVP2jQVN7VOuUiicTHRn
T5JDCD+ScvD1iEuMV8i8m9GzsVFuQ4rQ/N1ySG4TvKo0TTVa1NfWsZ9qpNUyGWZd2MYppIYWUekq
Mkgi25m2WuCZk2lXuRCIscwb0+1vz67yVpX0kDH/BfhWa62aTQ6VHtFQgw4AYomWSyw/Leg1zz8/
4o9CaVkJajwgO6QajjLOEa0L1YQiYgd9RFM1qgJF1ob/Ip/iZmZjCH9ZabXhkZyTFN0lUBEFvYyl
YPvTa0JjzIdW4mkrDTOJTRjoAb6HnJGPGcxXwk0jDK04olyMdsOdqr/1zDYaZb6KVbLce3t9L1Rt
LSKL/DD5VueJSfAGQh422U9kczt0NXPovPGyzjzMK/duK5tLJb9sjOc/Qm7630ABDl0Hlj6v4XqY
SUuyXTB8WHDRz9HtftCBrd9AMD7RIZoG/CBC798XFARrfNXLGPl9jpCld48913/Ys02LNYB2DiBK
lp3bEfbLEj9hsu156Ih8gaIMJ276D4icWR04U4tlFDFtUBbs8+AwDtO6uKk/KzgaWxY0e7+hJLAD
pPyg29AXNmeMMG10gsWzinnNSkOSs/1ud4u2cBDZ2f43VZ8tU2Iy/rtSFiAPhxmVr6ks+R2m7BPV
i/1U2fKtK/yFMwZULVpZY4J1NZXSWjXyone1pW9QZ2d/HrTFMOb/vA7lY9GZxVt5N2RMpDTi69w+
SiuMkxkVA34t+ajSJuz7MepiePso96/uef6Ubm6hc7olL7kH+Uu2h8kHKuyYH4N+MsVr4J+n1OgN
//yD16Bk+I7EHTHLHXcr+ygXkje/zBhwYA9YGHhTcOLwp7fers3M8a0VWfBQ1tfeJYYoPXDz80Ho
AlbBsXUBqy1HNbNZcq9b30wneEsV3qdqrjfAfIZEWclv1MPKV3X5MzhbtRhGQtCW1PzfpsbaWumc
3O+9A2AObC33dSfCPjO09gCRnD8149V/JPty0rxeukshV4TL4CwhipvYGfOD8qFpkvfPDadFk3bT
knRVhdA2t5Gk8BJwbqWSgW30aVQpfeXj5+clboePmadc1o8aHHceTZIHsoPtMHPM+eyIr45/9rL2
fnWxJrgJYt4povdvcZhUYxW1ooojg7wHOA8tEBnpcUHKrU8iQWCKzbCGwZhcD2ysCFBqWAyJmPnb
UbmznF6dCfYQq2fZtdl1JcIvTcNJs7smJxGl2d5o2FP+aI8hAXKsU/wch8DcXHYch5P5GPP2AouY
wZl6L26/gzXRGlfnJZIy/zm959Sgh0+TDHpJ9jW/AW1OqvTdRSgU1ClDio/jAw7IJUfmmT2EXnhY
3Qmivrf7ASvlKcYKb1uVgt96nQwF8yw8te2HHYAn8peyj2o7oPNfH0VqW4kOo6cKhymEq/0Hj6Rx
TLwRSm+bo8BvSiDPmGzGZf9pQd7heOPU0FHI/PEAj2N76j/TuFXDDMgLKiMlq1oxhBZNLQiBrz/b
qbZDBLBxfbyIUGSWStoYSapbPUcQSwDmLEY0DQNnFMVMcv3tPHYpVxycr3Xo/wEx5OVZfq10mmoX
6bRWheMZoVEzJw7t2RH17K2E1LWhwfvL+ePm1VfPEIjn2ujrFcCNgjze+62AJj8RM7cJw/am88Dd
iYUsisfpC0vemt/LEBsNHzION7dXZ2HCb95+HdnwmRSF/PpGL57s7M8lj8TrrAKlpTtiYFdbqIMQ
cdQmwQMFTcGJ7PIo5abKKZ+b2fbV9DtugDGAxltC7A0CTuvWVzbJ/Xw4G9AzlYHEA1gXRvzcyj0N
gwm608KOs5odhQvsuQ2iCCBPIkSNcToX1dfx1ihVN+22CVQWd/nd/ns3agUuXMWcjZV9Ee3bVzTK
TIUnM87WSsOawBShzzG8V7X4STkX7j8Xq72n1geWOdfcBTQJk6UYmZrHSagYFOxFtTuu3+vxyAl7
oOTb5CYji7QjNGciyYIfwpSbuDL+59KTcQ7xSRH7ANBg5sbASxm1dKjlXZOaTCcFIRxA+iS/fOdW
EMkGoAVh+VZtWuYRTLH97PDZUenoNZGlffQHRsqNmuze3gAbjyj/znJS1/DwifxWI/6jdBhjELzN
LKaivYYNbRG6fMh/P280zFl2rr+1D8y9LW3DOvy/BUHKBa1EvatJZkIlHPlMpR6LC4vr0jU/1KTq
iQGlsYYlkzl9hdypyA8XP/Bk23rR97Y1Voar9o4DYGjqkq2T/BnXVyR3zpcd2t09D5FkVf1u+q78
SFdM7LHXioCBxbbUPUvDvAI10IBp91d8H3DTSuHCJDB6MvM8qHT/1tfdGl3dC4cJeaTAz/5ztiUn
zasabgdyQA809cVxrJz6aCjctGj5mb9WkLkdin1cjywrjmMCXtNK/a+25F0LF9PdUo1pNZTjhqif
xEVybPUuol5OB3vLBxGRiKQLwB2o/eWuSxi8hi+VWLgtQMIRp2IqrU8mWVbq1Ptnr+CgJhwP7l+j
g6cEURyCxIqm61hMxIWo1OtjKwyM2F5OcxV6JG3nYCT9kT5MAoxqWVzri082MqOZ00f02as9zLm/
Xl1badMZLWT94/ZdSq0wf2KaSnQp+cN13KfqR3GgoF0eolWjsticokz1eREIFv6aLxEaJjQorOM6
mGwk3/MSx1nZAyhERIjjRJDeBVYJEhF0sxkrHH5C/KlFK6ZTlxheAl8A28JJ9NorgCYafoUnh6+E
pJfAwEigRMZYOvNWeySCj8+Atykclhw4XJlpGF7mjTkXB3jKoxqQ5s/pwCu00+B3d50Gjp8LrbXv
UO9V4n3D6fu9yujYbgGA67E6+Yk6BuVEoq62hl+zMrsuopdO84HeTngafYK+nLcNlNxMYmpDYjOz
F3iZOG7YJzdILU8vmMkb4uUEmrjxdDQD/TP4l3H7l6FHQALSwiwTNq/SHze6XM0nhAyglxH63vjs
7gUiWOipiUhdJNBLf0jOZ7MNRRgsvCfznCZvJ5pCTRML8bHYV6ST+E06wjQrfKRFsWx1QFlsJjzY
1a2mrIxsjy3w9VYBh3yU+f7kTlaFLgBlrOrpzV5FJ4CXr6vlFwgOnXwB2BiOvCeZwnRlw4+zSyWP
gy0pOHHA6wSgGtj7+c9M5NgjMoFWyhXi7E0nZkDrr7IG4P+piFaPSG8GEaJIsDfqmdLNPNsjkGyG
OWjQz59TkV/+vpe/YyQBHNzbdwbg7ImqnoJ/QNXwYDY/xx9SmnrnsklVJiYYK0e9lRQtWGaa4+GU
6h7w6ANQElOGbOgncjrvaY+iyfsQ1OmXcTK6/QaglNoykwPTUH/D+Jh4H4fbgwsaDoHnwk2hblmm
7M4v4uYZcAItcAILbKXQjmhaDIMD9Q4b/R9ZQZlxGrWSfUeR5LcQRd5zRT1YCZfzmp8l2uBCnaoB
VyHOIf8UMnl6ZzKwJPsSSrQ8GsT6fzQh0pBt+GUUFmkRpLk9si7+/r5DbRKEq+fnMcA+34zjCJED
893LWQaZJtKZiR5N+RDYoFlGcs/WnK/dKuCBGNzBLnkmFc/5JUE4Bd+LnAvH0T/eK4PPSJl0d+47
3WMzSAEylOFGZhTH4fqEJkBku/e7sGQyVf2iMcP2hqkmKVbZhj3A5OQnVPIQ80bfJPkj1trHJ38k
nANpD80SRa6DRBRXsFMpCzaqRnlG0JPFiYSXs0Chtv0uBb6Xe8svcesuiUhmabq4HnXIEXAnZka1
FNHwgj5/BonW1Pe4pPduz7whczb5tEBqQQ9ZMm+nlJA/x+BBLNrZStlHJPqr/VzJmigDySAJ4AGp
xSOVBSzYag3TsU+wzB0km22Drh9ZBMUKFfmRcz+LfDVATGxhtbwSVtO6J2HKZgiKgGRcfg6wJlla
X/dTgW7O8KpKIhE5MFeiktkYeS0JM29lTNu4M2ab8L4LjnJmxu2W6d2jQ7oZOLK+vuY7K5Wlh6Nf
uNYyWmvBkvVZQhKqA4VCw6D0s4KbmdPRM9+Z0KcKtKqYuxneaRTip35iqKmd/VZgLz9A3m/75zFg
8e/NwhTRAnzENI2K0NfEOVVAURR0jEDOnjJFEwpNh5Qpu0RJ3Am2GdePctMAq6PLRjL5ZozLIR+4
R2nCrUW8wO1FcyT/0mMoz7K7G75NODoIj78O6onf3wVAqzRmbr8aO/uIK+YdJqiuTXU8DtggJgqw
nMWuXEZPvmh+4LCGxhMCWTZl2QN29zfCDpbRu4V3P/J8oC8RxLYtG4tp8IDGO2kEP2N3BFi/eoFI
4fjtWAi/cF2ck4PNmQFXz/yeSfrliVUcIHBXgEalYSEaa8TG/PQj6Tu6TerJI7YB0iKdFKaZxJLf
x3neosQcoggUVD81gVYSkbP2DbCu0l8VYN+l/pQir6+pNepvR2b9R242iU7fiOntIrhLVFJQSTwT
trtvgIU5G8smEnXuAmJPz0cI8hO3QF/kqPnULLlTh+slcaVJn4ALORnPgUxTEELbVLXaagRiy7jS
5jsoQxcVCKGj+E1BBsNJqX8zUFL6Lpv2tSYg9cCrdM5brpk1AVvEbE5/fBCUhVvI1Ar8ABDPrOXv
3j9crRAkFcxESLD4bIvdOEkpYNZe86/6hz98YhGRhi05o2yyKYrIOGq0uYCb2EZogW9QsEKNMY5b
Odwfzyr0mVd18j6Pdey86Gv+XidlX8bkAs5FbKCEgALi/lMc+S6jlCdqoALBlv/FJqliqbt/texa
0vfGVcHapThwXR++Wvw+peaBdSwC1tFpJF5orCaItLhDXDQybX4zjKcfz4CHKC4Dd1B/IKsl+6rd
U2pQIEjhlt5hZXz3S5t4YBiUt3YccmlxLI4n9YBexetQGDz6DhpKkeH5KUZsAP+BPgDvQEAjOcTF
/emwqjIDxEelrBz6gDlNs1AGzyIC/lI6b6K0Z3bJLwCAfTzqkwI+DXONe/KGjSMJ71450cOUlcG5
008RpRsMCHwgrELdUbgfNL8l7qZpWQeLLSDNcfe0KIMR2e0Jv7XtPNHihUVKCnwgL83OYajjBcMN
89tjTrUw3kfAzKmJpF4BhrDiQLhfZvBO10Ax4hrdS3hdeAEIPBdRQh4T5jfew5KMCQ3iSbhov0va
C7LHGzbKIUzcBt/KTCXDQVdP9FTO7jXE2mx97AxMStBQgSz42rAkDGq2FhokYixP5rn0s23d59CZ
McYK21WrgncT+43g/5xDSiI7ofLLvinz2gnRZkwLgeIAm9OKPu685JQHV+pT64pnvZLcQxtMVbqV
cnIVvQr7VLatGqmB8cixA1++vQF3ZKDZx4xIXHctHiNnYKatv9A14vQIhJy7LN3loon7USwWq4pZ
Utgav5IqXuCpCryVXND3/hbs2Sh88m1NrI3cn17HzSc9EGYg/aUV0lgzmr+OTsQUpXFJH9HurPAp
/LVF3JHxaPrro7OLJRr3STRvwHssRrEWwVP8WVIAIF/RIJ89HrBZ1m4WwIX7eUmYFsYstrf/26rh
Sog+m/Lg7+jBVJ/g48zNXEGtRzS0HerZo+cmolDkjD7IlWTJeQhJLMFk63lgqic+jDHQOMvyXffO
KPiwStfZ6zSTkmF/hJKEDrr+Yhxx6u42ZIgK3zteiz+Rtv3FFTm8Ga+bvJ7L8uUIhGF5iXqBXKOn
bE28FAYQhVGcjczlz/mV0bf3HyZhsRS7paFCNDzKnOKTsV50eAr55NgBRQK9CPgDHo/jpYS2wVaT
V4M0fdMW7a7hXHcK2uIhwl1tam4DJStYPkq6o+KdPxojIhOZnPBCEwFWb2klZaV3GsQ/zdAccJDZ
wTB4uJLXQoulqvPOEosXhhquXAfYBVJgwOV0upNXyFR5m9+30l1wqXOLBOajma09fmaqgsX9arF3
YyOYGCLbqAT/Ga/UdJaI/kAgCNxvJNCbPQ+CPMmTOLhXrvpusW4IW9zD2VfKioUqU1prHKDca4q9
uL/5IXWaD8kuQJB/IGQfdsCzmTNH3tk6PQBFBLqafxOd9mUWy9wZvYB7jgvlFp9AsJFbnyywwI+7
roRUs/m6hWYOTwUH0T/Wxv5nvB7NPt+4LicKlUeWrNZPQu5uVb6zYqAcXrD2Ajiq82iTWi1mXNzW
mbsK6W/BMOaBFt/WAzJiSqW1IOt1Zuo9BCubm96R/NQyB6jTFFSLJV7xykTdhWEAitm0Gfz4h/Np
mT22fNHTEzocxfsIU6mfebuzqoK182yQRDMR9wVmBgOzHNJ1knKfx1cn20smRBmCV81YXvDXf0kZ
RHpqxKkwI/JFoSE+Pp0fkOvN0stOJKlvnpE936rcsw4QZscdVvq6WQdVEKMtU1Z1DKykcp1OZNLo
hk52d5TAPc6RUvIfTOg4Xe48P+VR9Yw1iW9bTj/gztYoQZXbk6NMVm4uxKpU15iQ4Mus5gp/GA71
Sh3iXNUBDjpD/CCMVc/akRK5zpI6djRdDlyB0NelVY/oPPpUpruKYjl4AgJTUe0fJOLP/Zn/dSs7
yJfT4oU4lpmxZF+FKKoU9HEKJ/o7Ldc4jv3QRHeSTcDeJgsssXzngEeezjyATH96a6PeSkFT6QlI
RqlWZwSAra170Q+isSN2SYzPvTkG5yvwwMqeCx20sR0JRiMfRqL195cxsbY0QifTXh/WDlCZ4Xjv
WDXmwujK0UHIdRKpLuENmLstadyAYrB3Zyi5TssEPzxJ0NrsluUEFW6X9eZh+F2z51Qp9HtMLwP0
sxOTG9IXnMz7k8n4HGJEleLtn9mkYaCkXGAk5O+cXY9EG4+/7lerz31IW5Ist3hfbwnfxAgybBDa
VXGJQ9UcQdiKZRrHN2IvNMvM3JSt27RuAy8fPJo3vxw0Oz4+vCcjT94Os2i/hmGVcdDSKHtD74aU
4xFb3jcwAj8msf4KrdFmhQDO5mfdZ1iyC0S5OtZHLduEUSIIK540TiV/prbHPOCfbQodlaSCKBB9
25daMVGJat4Zff4blvoQqpzuFwNrNNxzDzPJZyNrVbOugpTCZ1Ofsg49rjOdl5qFxcdKhTLCxZl1
zTVuLNNfJ9pdkYPIZSld3ol640q5seU30Ui1Z9cGskbBxaR6GiS/S0bmu9iHeMJ8FMNX5rK3ovWC
Wgauq1WyQkleCg7d7vT1/BzpyoBJXHLkawAL+K7PwD/jwBQBIRLmVs7KrDAfefQGyJMCG53p6maA
N+kxWNUV8fKg/ort3oZ3rrLwPc0XcoLbALBN1iN5WDW4VK4ScMpMYp0DcbhHmsrxf3xcSYi8tQ9a
brhbHoqVquHvgMKTwBbWJ0LsEtBg2StX7K44aJVbtwQO7V4t1aoDry42i7mpNjqgvQ+y1TpRLk8y
jXSey3VEkbejf7x321AduT8KCYxFaCxK2IhbTXNekRgjbi85+KhO/kY55gycin1a1hYnrRRzYtLV
ZiOroRQsANbelJQOlm0fgYTXpt2al4jB1Pk+dn5pEEroWIWwblCnYc6CIHonLOSL+Ey5EFIHYU7S
XJO8VSI77gt8S+H+HmcKuOmBNHvO9OEOaFFAhbBdFdf0LENlsYsqVUk+ZdSClYS0FEFhDq/LktF+
jjI3lI2T8GfTu+n9MVsQkhNOhMtlRkcLwEhQd9q5f27lm5fQDARYX7d+QS6KFh86SR5RnKE58TMv
cBB98U7hJIh1OJ5DWZ7zEKhm4Xy14qzTQaN4gGYcYMxXCnOuAQTCr4NPdrGzSKGGOK2SDgrCYwf1
nuUrs+t36RBr6oGrDrEMYMjDwLAi7VZz2QAsjQDQ4AWEvHybAjELkOFRc69DYzzizS3HI5LdE7QC
kwYK+mavX67pApeXErnyyT3UY0SMoGFsHgXySubJomJJ/WOyk1n6ItM8RNq6xAtcBqopGOGZo/yH
10Bkm16op/mOjd3cT9mykHGbQgKyLXyPIRAx3JkxeBsm5guKzqlw+q0tlIa2iBNvqwOsbH58rPS2
YXa/U+8ht6mnCuCAB0QEyCUXVar2I+QAScSvxUSXujP9JvmnJpp5R2+Qgj+xE7P/V3o4ldBk+TCC
Z7g+RxXvC6KvYJ26aLwlo7vhf2LPsFva1d+hZ/xv4sSEpXMK1ZiWGU1L5HQSeQnEEdBggxagOmBC
H11mVsNRFdorHN+bjyt4q2WOT+trjkT+l8rXHkrsquM4FhKeuO5vTz+PZafJFu5UGZJOHFyZK5Xd
ZoF8/9UQQJjT7AU4uc/uvw0sfwKYlAjELGcrykdy4tTumy6+lqZ87xr/8z6+lGi29kUUNdpby+XP
CzGuO3Bd0mOvEbV9wMC6TO61WMmdR8rcxlNhVmb4vdK7J1g9kdMaRikumAFR3zEob3BUliZXlJVu
b+HtFUDs5pNAE5NYUGKyyF2yz3RRubXItRYV+qbKut/M1snGRn9OrmppKkpGFYnPCN/vOGm3Ns+s
wbtt0ZzXfv9z//WFZz4Nsrod09mEo9bsflLaoMArO5m8uggImkurcwap3KOB8Ty73O9Qq6zXO/5Y
Wk2ERfoyw7uGidKInJZAaG1gU09uo3dAqB3h/mnek1AMsjbm4kpJirvZp+fgjjQ0QnQwGMrWSzqE
ULsY89KknOudpiMgJfBpwFLTeJ0mNU0PgvU2sL1IWf0mOIU15Cq+uyRlsXvtJxOgxGEw59zbWyZf
AqhcDbufKcVxKXN/kOy7gX2HCYktHRfp92MDw2K+ythtfCr7916BsXB2QJSKlx3uufWPUOmRg5Y/
XSvSxBUVfyEjps/TKKks9iytlB01viTKIsBkgTrlPVtIlHxldqHnOXu9r0teOGXZEp8s6dQRsTiI
idesPBpCxJMAmiVlySFuJmDjbLxasN8dfq/KUCV/I2HUm7Ld7FZU+lfHjaL6PSNFxsLpgdkyNmJu
2AAxToiZGj4uRu6o2HqF2nBHogMqcZ3XX0SzxSu8bgTcPTykCZS0o/6DhUkNcP3UNs+627+hmsL9
nwpdQQkbk7v0tBjHUN3UQ7BI0C++MTtdBuGCGWBQIarmTH7tig6Wu3pzoZwOPxYZjqlb9AMIN8t5
7yf5jnd7StB9QP6ziizxOOah4QX5ZtQoJr7k/3BOY44hax3vhvi0dTIsQFqhXeqPh0ewn8pneub0
cs8jYfeLNYjlmv6AsNptLlRVcYVqXRCxc6GPYnn+nHo6UR98+LqXkUu6x4iDI3tjN0dyRd6dZQKC
72BNZ+v3wmNve+hnKXtaHH0hwBLsjcc+7KeX1X/Q6sPlMQU64pnkuwWXAfQ+OD0JkyX+1h6OY7uU
E09yiLhYgm4PQuh20sknAWEGALZxhlh5Acv2AgLUWMVX+R9EMQHA46Hi/QAZXIa7niaz0er5Zfrr
O2HssEABk8wWvyJXb9ayhP7O0iQ/bprCbkrIS+HcQ7SN6YyV7EORafWSIXxkZMVpTYkPHCvn9o5n
NqZ1vpVIp7LdkP6XSlOuSDn0gyZZuYICfnvYOBNBOPjMLJp6au+eYfoffJxMfnljPttpop3aCxsl
R1sGGKT3kJSW1WHzj6bxPemDqZHR2v3CEKaUTwg0ZlDw9Tng5kdj9PWZhEeXGk76Cs0eHvhJhmBj
okphVUU5oSgMjsMfoP06Ow0U/QZuf6KZ972LGWc8jJhhPsGLDHx0fF1cDxk4NTA3wc/Ir0YqSKHE
v11Hids7NUkc5JNR5uCiUGqUXd1auFxNI4dDibHKTm1qlFtqT1jMd2iNl0zg6O1kAv0YeHP6vEDa
wiJl9K/6Ir7BL00ffHYsPhdNu1anY0MyuERHSeFVWAHKtm5uMDSZDRE8ghurP4qkoguYhm7/RooC
H7Gql6pu10spjTDXe973h/6pJLFUNQuld/FIaPgEAsar66FLyvF4o5vz9cu6j+DxRpDRSXSd+upi
MDejRcrLzkgY4/xAU7zZlR8tXL/7uDS5iUn25Be3uxNhZdTxOWmUTwxqy9ULzKWRBmQ/r8Ak+xcY
6Y3W8/pq/2hSeQo+h9D8hd6CxNu9FrWp8LYGIrZuq1gYigO7i9hfiV2X81aF/mf1V3wS2vpRZzrs
1X2gOm0wOY2pNzDELGFo0+C3eJcCR3B8M0+XAJH3FMwCs2P4Rg/Ep2y2+0uQPr7I9X95+8y6xsSt
VyZm/S4JkkmVf3ZvUZDp2enkz2u2k74BJRt/wLLKWgre8YVOX2FZxozPUM/ZyxeI4Bn7aONFZPUU
I7QnwOHZvi15zh2+EbxvKVlVEzm1JPYloXze3l7EBFlwWDgIHWSXWogXhWqww7Sarxkdgr4iXxP+
yCx3KyPIjmRgvqG47a3mvDgyXuIoR/QkLCPvQBdjLqB5TEa6reQtt0w2aX57MO6vhUpoRmkM2LPr
KbzW+H8D4cY9LTvocDG0yxqzQEIHBZfAVuT5QEKTAbMNY7CR3H/tlHAVsqHGBLZ1nZYMKe44jiiW
eNoku4LRnXlftkctylhs724EDxKMMtBjQvczj9a4snqIx20BgJmqR6FbQvA8VKxG/YKPk/P6CfY7
LHYFno6ZN89EmbK/HjA8S6p3y9PY4xGiyNSoRYk0ceYYk1N5XquosGNRizv/WM1hjjtfqirfERgj
Oby6ZuwDcMwbmSHfLEaOSGXlo1D6rYJxKg96kKx6U5YGj+mTP5nqAmmNM43zAJX5hXRKVuJFg9vs
08nQveq/r3z/K/eskc8uC1nOjX/sOEaYrq4ck4m3iOtnUN30MSbvHoW/6MSLFjN0r6Ymf8fUmNkc
dxIqMeVYkMxssTwz16GGHZRXTIimWBBJAOZkYYLP/iNgcMV5f6wDAw7vYd+AZZdNGs87QLY0mYhJ
gGD5xcbOTnxu5ffSZ9r+qIgoWy0Bt/i9G3qLvcmZP5pJ2Ad4C46EqwHzo8hmBwi2Bb5lUPOQMs10
KBWa3TdzJDbZiaI8H1Mpuy6zoHWBebMhgMmPEdi7TCrIXhiNothDDkxn3S6BIIUTmazwIapGVdW0
4IA92OstlXAYJ4xjZwGwvDSmSSYXNj0GwrNE05DGy3eGWjtT0l6BsVhAndYZK2E/PWK2GR6GcKJx
iWuVbvu/OZAHAro/ht+paolreEXmNKStuP2ZORHeYZ08QFdy6+vrd5RGz8RS/fHQZPGByD4jp00Y
DHKtgvjfVatDiiXGNHRjrNbJzLfloQ8wvGdqnSST3dQogAgKO+GB5pIBFgpowjyqHe+NDl5gz6G6
n6KfP0CtPNGNKo0/ogjTAl+1nKkP/8YHM0g6Mz2eXmt5EioxWTdPSQrRovjiNd4BBfCuGRzrIQDs
D6x4wfTMuNEYEz42SuaRZIHpaddPgyuYZOpalr/6o4COjH+I8RUzXp5ZdH3mow3a7hnu9nfMa0kL
Y+oTFcyLcqqxf37Vpg3CLHyDKIGXcTxS+illnZKaSrGYTGpgymTHwQtNYySfZEVunNQ9X9od9N/4
eb2zsXqN0clBeilGCbn72MMwaDWbg8Ms8/BbXd+km8ajLvbGqUiBIrAhlc2vonR0HlXxkb40c4uz
jGBg/FLKkS9Fzc03/u2iit3OPQ77iSfCUcglwr4MzE9MC4+/CqZTNx7/yunAYUJSssogKUk7Rq3D
2kBAGEaVB29EJTtppiKBoUqnGoltAvN+E9WkHwJUvyeYW18Nki2wGfJKwldAl+ojI/WsR6OHJbUm
vyTpjo1yHQu/H0fOmBttDZEFxdjkIV5kT8JMFmigs9GU4sa10G95oJd2oYgrn+DzYgdxVI4cC2Fp
PLYQPAMp877CedGHvNEfPFwHYwsfhQFWkrlzEdlaFq6B/k4Sg8IZ5UVffubkFinqVq0s7hr5DYT4
yyhnN6j0kkXdR0fmnM9c8pamVikdydAb5PD8xGGHB8NPRndnouZI5ZJayYPPbvQdqAX39t2NLI+y
vriKLbDdOPXBctg/LSveJ2lnSTd+JgQ2cndWARWs7TEc4KK6u98Qsi681Yjh+qEwYTGEuTVIl3ub
pTZCZTupUoh9eVULiYlATPtltUa+egRrfntVIbemBBzh9JOvKo0owf1fxtc20wE8repFFMpKb2uV
M2foLICBdU8TjUZnmy9C4myLX8RwSDzniR2JO9KW7MwMDvG2M79Z534gw8RzQCa7p198+wrW9gKD
x+QtISoyOCk94WI+VUkg7TWDWITQz9RV2n6B323X1JuSPnfo+hJnycy0k+cMHCXyWy77isfCbeNT
Y7kQrhiOvzLmV3ontplFncWhxe7XmI5XwmMhhFe4TysII17KH/PJCcTwG/rRFv39xvPBaj8pxNer
RcXMNR6C8r+s56ueUqvM4p5ZdhF29fWNQGM7M1KvWmM+uY9PsTE+CbTF08MnrblH3j3UV0JqkAGh
D8VFAGF/0waeq7Kyaf9OKL+EUuNKrTCS5psH0lj94dm2hYcQYxxOfIk8ApXiqIomaM0o3b34kzTt
W5lk31bYrrvMblMekxMg54vybl6krdDEWk44Ue8DjDM/UCjDoTCDw8vP9vwP0D8xNlP4VhlpRnRm
UgeUwaYAGln9sDb0ecOp6yF7jgJNaA66MRwZ7W5IN8qnCxwYj+j/A+IhC0izLDX9HxKDcw3Wcxbw
gnYyT2GMgpA9wOiPUCs/mYdm8jxr7xrYh410zgtb9MlUkwXnqbC5FHxwkhgFvCgsFrOcQppVTK7z
uiQwFAbFApE4zVaZXt36ag62jks/qR4wtpKTMlBjYVYrLXPXiAvRJ2LwGnWNMgGbIJdNEkDS3ciM
aok4+8ZaFk6kd+2lyim0QOwcmCYwvvPKsDCqJmcegEbSHlT3lNY1FagfoQZKQn5fgjN12cm06Yli
MDRge9iAKsEZ2jp3jRhAQDClstWxJFDRaKzFXkg5NbvVxwWTGnfaTGhCtyv9ouIpVJ3RygtA5NiV
kWJxA+L2vGqE3AL23O1YEeGazYpjDSRX+aSDEddMMpJ4deKB9/KSB160GquycIJKJ9pn8UM4SMTE
jtrA4Xj1+hrRvsVgSeNPtd+PA9cUl6lRJt09xxR8tZC9xUUT/+wcJRjF/yinTB1iDXEbUPLak04q
XRBZLVHkwmB/DkzyG2Nzxoo3PWBp2U9842NUGZ1hPJ8+wWSS6BSEnlTVnHv0p4zo69RBDUrzv4D9
5p7KxIf0iMyhgEvRhBiUVreuFaM4IHcM2IJLIKGNIxtpmEPqJ+/iTtXM9qzMyliRDDsua/Kh+cDv
Udj1oILnRUF1vzQDcHdJ4VoSKBZqRZNGbyRefsaoYmeseqIVafZnuUusrSNXafdac3RgCQR0khb5
Mvnq+TSElW+glRI8o35yuw9t0jXFPoJdVbo7+vWojDrPy863+WRrn9lYllHu2h2q9zi3/tcrKRi5
aBjPkpsjbpJ3CPH8qX8NWYrcxGc0xVW9u6g/Z0x/WhhW5ei4L/cSbswkzwXvw9jtxOjj8x2yHSJP
x0xedkG+Exl/IhlVPQN6xX/n4X0ipD4EZen9xV8xjWM0TAyecbskqarNEpNnPolAA8N9HaPIrbxK
X7yR20ZY9FkiYTsboMFBpIEaJCf2T+ccDmaRhLkZSS+5YpQP/4tvjFqLKaCkeSRNx9BsdbGcLrA4
muuheR4dJvXHuULo5AIvFJjdcvz06QekFrDFkREFxnsio+yOIs8f5mSOukIcW8wIqUPUex8Gb3NY
Zu+hftWgN6aczFmj50A0KBoaf1SC2QvzBYkADRT8w5fxPeqLwiFvxogj3SzqjAUz5JDkKVnb8uqi
ATh61hIqWzOilTaUlu4CmNB7TBlFM2r96MzJ5gJwDwqfiMWctgn86snaGWtzGGsmA5ZkAYtOLY1J
EXxRuBO3Dqb9SWtY9bea0Aj9W2ZYIom6AO81yr5hVZy2pnqIpfTr8q3qviDcRtTYL4/lQl46I6u5
bVXnWp4RIqdtwoWKmLw1F8NCKjuyCZg5vgM1i6p96QnSX8wRMqL6tv77rm0I+t6bieBZbGZavYJX
1JEaVKlbwsYf4z+GMfjyZoeBfVdTeEl5Obw+uoWRICpDdmNPWC/wz2QspS82Cer78S+RxLlkl0bY
XYlEN5SLWokDPTEdwPJwJFc5wBAD+8c4l+aqnvw37PHDW8iENWJA4sdRq6IZbhmt+0K0G4qDC/8S
I2Z0a3yPW5UcimTs8tm/Re/GHx0TN31D3wwGkJCeezTUI/c/vUNGQ4RAfJ3j+JPouOtubCQfuC95
6+5o/LiQv26Mjpv/hIeD6T6Y9fr7Lk82V58yYxgNAIWsaItW8QR+s7d0aNBLKqS9Fdm/X/WZG0hv
1bwSbiEyf3UtfZdtugpB6zlMtvwu4W4R1GTerOSfN8UawDdyp8CC8C1CcfP4FxejMOVpsUSoRiAI
cxYUBrUDmWRawOGptZcMeVhaWjSlACPlKNFwvGgzlpgoGS9yrp1sQ0y/ASRoe0oYb5M9uLXlaw6m
Wv5kV04t4gTV6MLaekZ4qlp6G8z58G/BL/t4H6IVetAdAPYoWYy5ZE0T3YDUC4gnYzN5RcUoEduf
jlfVRV5VTEuRqfT8ILfvdd2Nqrm2aTsaWds45AhyC6PAtgRL7P/+PxSjlSeddRNQ5UchoC+TsDNZ
f94cRtwSo4vKQ01IpLnYJvxYkDM3GoqIjbTExsnEhNRB91M/PCmL8N3GFjOk5NsAzPQU3bespvWc
2/mu32+92VX/g+7tRfV7P019ixup0CXc3r7d66aR0C26iqo9uCR+eKsMJJ+TldwVIaYN6oWKmeg+
xdspJ/5UwZl5rAfffDUUsW4kHUmkwF0JfKyAJI8lwiBMQeHkmUj7VBPG5xHxtM2Se81GeSyPZRE6
nBEgZkKjLZ6CW1hk+an92oeqiKrYKEKV4hnXszcx9N3PZw9WIJE5+NWsu0KruvTQrgFqWtd26SM0
HHEIQPwvnh5CekPZ7QiKVBwagsH73es8KG0JC+UJKEGeb+U1ZWN9a5QE3Q4HwrmGCyD3eJudbfrm
YmqL6jAvMIs2hD2FPrRF0czeGM1hEzOV57eT9h0yN3fDNLFFCv4fnvgrriIrv7kpbLpulg72+Sie
o1d7a/e55piz7Um0Sb2k3AwMTO1KPvXBK7aiRW70waxng9sD4B4nyjA/J8F3cwJSny1cL5DhDQSy
L2aly9OKZPeWWOv9Zp71Nwh3uV7QX80gx4fMlD9ZDvvJiqyAP1uOKRLvUia7W79+MCl4GQAIUZVs
dr4JDNwA09A5RGl7JMUoD2xVlzQv0kU4hPKzs09NdLUAVxXHVSXXgoCMItCTVcHoAMrlM7b1SH4W
aJaZ2SV0n6WCIm8Hq9N+c2Cka2CzwXfNWvCPJgWE0YXEvoJxnu9dtle1OVESVNtO/rLgBq1ht3Jj
EHVDI9s3qs4EMPolBw5f/vbM/FCYv52he58sez55nk6Io1CW3qzWLlxFX9yh80pYjD0RYVOD3p2e
BVwDDGMKZgSrtP0PmER6Gqvj9WjXbqcFffNKM4yaP5K7bduOBbJg1j4wQc4RnqMPmturoyzmAP1J
Pp7ZvwsT4tFlA36MX8Bc7KzxVpmweW5vEph9Tv5GihFCOmamscxtY8k1GhgpdgK50jS7zDalgRiA
Ze8K/VrEsWB3sTE+Rg4kWlDkOx6mecU1wJkage+JSBdLYBzIK6/1BqUnKFV+b0ESdWKMl2/iSjuy
IsqgSJxHuH5aawzmtdHw69Wdx1qPDfemH2KPrVnCs3/BCsrqm6gH1jQ6UyHp4NoMaKdXlK259xlR
QNy99/LM9kJultWV5yCO9d8dEi8VljEIVPLnJ4sIwPpi+HyA/yy1f3zaCedjdwoF0kFYrXm7mPhY
fGhC320Lgvxc5Iv013bzsseWPsH2ugBrD1n54HcqPG565ZDFkcuSqSPDUMIj6y8F2Kq/3dkUIkDb
y3RCuu2RHSX8q3DmwQoQ+uRG393hZezOCxVAm323r0BdZc0sSPXM9/vg5/gRg+DCCHBVuQfEsvZt
2DXP2VL0BOhjOBm8Fm639eUzvB+yyH/7rXTtGx+NI6K5AcGGsqUyr6puTrkwFfPx6AGVVyv95/4i
oA1ML35kZxwYuho1kGNH7djwSFKviDwy9HVtCgPAEQhP+HwtjzFWPuVHXE4rXVLHi7+AsdCrLNkf
RFeTi7fTHTD8e53hBw5sgwtriZmaG+LAh4wM6rise+MH+fNEsuku2qsGoF+taSaA/2s0HjSKlDfb
i3GwiC05bUqQdFuC/n/zyHJY8AwbzvULaQTzak+kgkvIeiSZhywHHUW0N7EnkkF7OPd3FZbCHmY+
WQbrbDx7fFcii6/YV26DhsPtF9zSLKHUNJxKDupNF/tNOS0ljFnklqQqY5KQrvWABUj5IE6jyzlW
UZZGuYI61RGGYYyPrpyxJ3x/1lNaYs7nKsjV1n4cZaSgd9Rh0QnEoWD7B+jcYwlTheVcQBR63+xk
XzCi2kpo6Vdm0SlNG80BMAM8eLlnTFuRUWD5r1EnjvnMDjCxbTq02rD3hPj+qNoa3Gs7V4pgpjE8
2kzsuxWGUzo5aYGeuFK3tGfF+79JyZhpiDLihYIy8SpaOGERkFbA648xQV3Mk81ymLSQJI+8W+4I
zAHqUiM2BgVMOgjx6xTVoRQr0VrgE/+Q2/mBIfqkJd3bsiKGWSBQ/aEt/APArd5qI45H7oaWMjvS
stGSe5TvG4S78ZlUt+yRREoI9xFlAHD7MPeMYOo7HER4uAj81A1U6Yoord/19dZrbZSHKtEsVjRL
6syQROWkdf5L4uYdOCpPwSMPqQntZa/Wftt9me4J0jonXlokKWzCCbhJBw5DEFXJRvJ6KbEMBoU7
sNpB/H09b9KTeotAszjwl86lIBZhfyJ3c6GOKAEsud/nvZOjn/n7bJTKgiFdZVC5hd4eZIVAlGsk
22G8j8GJY+yUvf9+C4B5SA9Ruw7HoXybhioNefnRsws6RNpUD7gqbpwdTXwyfpzPny4bix/Ae8vd
p9GZXkdWW82hueSHIUZtCwEj1IKtqysSkRb0W1SSol9x04ngVgbU/TVeuhHfPEONtSiLtuuG3r5x
jvUjCNZ12rSago7tYAdEGCEFkdyio+CFIRX0dhH1jjG3jZON9FkfW2sml3JNJJhnn6SNhjjGZlSO
wg/7FVjt1r4KbdTPQEFYs/vTdMd1Pyo42ENGoQedLCi/KNdOr2Amhz/npr/RqP+WXas8WPjEh+yo
CpXnE7XAyH6+Tktnmv58HRv/XMLm50D3ezK6Jlt4uFBJNAt/mkHo0xTkoyTHzMLXtf/eD+NJKIIz
3MNyMMfOGHqEhI/b9prLRPrBOYe8i+sajUr0P2Hesmu1W4ymLyORs5dAGMkwILrJ4D1Wg911o/zd
dQVeRe7Tq72kOvdfBz/33Fmgy4f33vLhoAhjSZwsPf7kY5Ipj5CIxCflALIeslxFiLPsQHl3EWW9
wXKe/Wraxy8uQDr97iecaatkH5l+hXBujNS7mV4zLNCwEhOLYSbAZR32aAYhTZzMslEtsbM/7Ise
vIvDQAoIrzZB0UxXfETyNAobUXUhKVmRTzKGdAmfWUh8QKqBvflfr/N9HgNdPmumMhtr0F6VuAuu
C8wgZ9Vkhh8ADVZN/SB3L7U5C+fc9wdcc4P74tV/XjcuQyK7a2uWZvNGlZHU6qlrzgEvfVP3+gU3
tIM20KAc/1n2+zcqyQm8gbtsnqjQClzNOS5SXZyMk3/CZVjljje9RrpaOkn2DvpHLK348em1LWGW
+B/t5E7nGQlgvHHrAxkZayoFA1nmq62RVkVedtmo2iDyr0+aTO4rL2TKTt2v2kKHkaRM1cvh2yJQ
zOUOkrErcWJ8DXXR6xd/3LuGKh5x3e/7/imyq6qH9mQIqMLuHRZh9DTbx3TJMBgqtMddcM3ptiRC
05HHV9KhEcPzMeRO6r9oBH+XyEfvNJdpaqhga4Vtvf8HAcZVGmk2fDoqfUCm7I3Wow8Gl0/IpHVi
+YyFgfpeaoIbsqRnyQbsoE38ZdilDbqNH1f2U/X9kmeVH2NDOpqb5gYDz4jyhMX8NBHzDNOvn/y3
BXHPhZW6njdwpacRx0O6e4ZfYCf4c5JTx0qTwKh2CwZPSDSYVQ1v5uqeAuE94aJt+Ym9r3NQ19/x
EY7lVtdIazTh4TPAvusn0zRmEWC/W+3u1W7Fb2vMYIi6xhzFJVW2N5ymdJWVXaZIw6bDISkTYY19
ke6DRkyQK+LVKK20pqfyUpTgpIXjNi06B6LFOurRNxibqyk7YsXUp3V8lXId7H0PZJcT4nmf9mNi
5027iDViIff9lboo8ywGORiHPb07cQWMQZT1eY63VxzW378VzSJep4TLzzoi4edvDWIYfBTU6be5
YHuOCdKdSYucjfNRjepb1LYnaDe/A4A8rFZbvHvubn0NCKHQ7Gbk1z0bYKmKIosi+ZtY1F4Zakki
NZy7uO+Iv1zIyJq5rmDuSZvp9I1X8/pX2OQnl/SkH4NMIM5OYk2L4GzVawfZ3Q3/TLLBl7ec3Ttc
87pcWyxWUPCk0cgmf67YuRwh1Z77L/uw3KzPIXNrJxWriyjVAx/tHlkw58tMWaKMNY4bDKEXy1Ta
BYvrp0IuDZnVXa0snwilV1BVtg1ePhbTq5ivcY3UdxUGGtB3Op78+zAFZW4EZTHQJFlZE4EkybYK
LcXNW86ld9UCJo1F6d79znxlvrtZmWhfDOSGppwzbakC6E0IaG0l7dwm9M/HiBJ3oLIHCp8rJ31s
Stt1DMTpZdXIA1p+wlpWjxE0QvcbtucmneGQexbDtgqAaKcKByGvjcNvAYPORiqcrrpxjAckDvud
ck5ep3bx2YrHeKFMNTPX1swGoaDpHhhJjglA4CmDLWq7Gnie3wwjOZeziuAz5TE+VL7uz4HlJdcS
m6U9VZqjzSmKIefFQLRBrukAr8rg/CgNtbPDAUBLqZXzrnuj4+4g50xylHlXePw9NOX5gSqGPjQZ
C/Hu3VRwX1wCHEp5bzIxB0hsNETVNIDNsUzJSh/AAY/ARfQQRVEASv/smxGUvGoQhz19Q26x4amo
a6WJyvmGCcS3FH64UP/zJljYqI/7l3Qc+MHyTsJyExComjzSkUfxj9LphPcg09jbiGgVUrJ8SG31
7VA5WFgtGfRu2GxnldiKRO1fyzwgLiLcJHzCi0Qvtxs92ssaC+LbuaQRsmEzsjNHQLOQpHjKm/pp
Qe8xV0TKvcTr0lI5k1KywVMwSIUxy6RztofKHqoitg5kSAHJeFvDkTUbCIGV0opta65bmPPRT48H
SC0ynMPoZ3+DUJS9AawiT8IGr9KuCtO1g8AYR0YNB9a3palmRESgehE9Nfm+71JzC5S9RDmGU8dr
Iz83FBkeqo33TBmc4+oJzi029LRqy0vPlTYdLrUdqnDD/rGWZELYBT1Gm4F3QYvrQRccHFjX2RVC
2C1UDrOv8trSsMRqNEHNotr2JxxLUjFqshWYQ8fQaZhxoa4aB301SNnhigpKL4RnLwG6UL80mrWU
CD/fpG2RNcEW3JaRGs8h9Y4Sh3gucIwRW2VZzZbSRQpP/KcTkCNiutmV3Zu9WSjtXiOWyCoZDxVY
HSBuwu+fTnKkO6go3cuFv/O07YBSb2VnTr3+XTluEeM/A4KYY7lF7nFYrqCAmce5F+gg3n6rpmtO
zQnKNYkARaFcPqthIR9oD9ge+qHTkir1ZohUeBjdoPOyws48apyStr2n/aSfZi//rETQPXklDE46
0Y4LqUhj2dVSZ9CH8MQ94CKcx0smOg3YXPRnK8mkREzhsgQ5JMcE91qts+7Q+2N8QQ0gArHZxDrt
xPn3RmAHC1oRKHYWD9V0iWPvMCYgghhF68cMV3v3ldACecBZAX0ap/foPsgjJZsnqvIQaosIuak0
8MVE2DKk1td/sebnXn2PkIQEvMnKe6t2mP6dDJHijkPQ/CLfXscex/aB8xc40fgeLumny9XKALCa
YET52QHPzbsUqtyoXjomSv+gJrdvRkluiCgJ7oMwZ/0LR/44g2WfsoAITXIoCVrMAvIcLSz7hven
MuIkAZM3VXdamBJRipdqMFnKCPsKsAZ7mPCMv1TIO92Cd0MIWnG5R2VvSNlf4yiGqV6Fnhu86kUp
+6Pa47WYL1pRBRj9SOldD2ffjd50tUKuYOEeA9x1YuTwnO+uSkRdf9Nzq7ImtmN7u9vCeAUCahGC
xMaIr5M6AmqoW4MkjjI3wID5Mpd6jRg3Sw6sSBlGHPGPm2x3WWR2L7+IJQuvfaLhPoH42HaakLAj
haOPNnnPQKWloa2UlKqb4Gqc7OxmpWlUFkwAc748A4Nqsp3zcv87F0I2bd01dVcIJ5MxWcdkGAIQ
iHY7hb8DlSPP2Eq2Du7s3IsR1oRucOxZGKwycnMU+qLhkoLvEGPA4j3yraICmL8dddlPvH7Byo38
jF1ud5suwI4bgSHveva0FxEcxvg3yeMjxJUAWeqqIqm3L/CSt57EMyAz0RX95INlfoGkAIl/xQCg
faTutvjYm64zVPDkv2BUk+VmqP+I/Wx4sgGJT10opUlVki97PT8Ngx/dCShwRRu/1+S08CejPQRy
QtBqcxboN229xE/8ZyLixHs9LP0Q9OFPQxkPeRDsJd1TfXwkqnPj38SfTFrvxSmlf1Cr4IRbk5Jk
T/VsSTuotNoRzaKmnFr9g+kfv0pGKqgvHrvMi6qRmRUdw75DenS/fE3DDt+Y3yNg1Hg1ank6Bs8+
AG/DPNdifo0Wr4brxNgeQK4fjfA81MoWeno6OWZfE82PqcbOFjxukkUz4wVCu87Lu0COokmUUlac
+FcPRSeeXn1GYpQEdgWnLcELFW5JBymVlDx11gm5dLCQrndx7f4iIH0oOsjEP3OnpCqLNumOMtWA
S9GlYw6V95XErJLVmc7kyPVLEx4P/F2GhF0rB/8XC9orx9O8m57gPHpVLiOZ68NcDqbW9C4qg6fT
Gb8bCPW8y3XYan+zmVIkNQ4qerXc4LxZdCaC1BaGkxsKsv1Lhs4WTBJB/akTorTtzvSdfJI3bXyl
tJYYejTMlKPMRIePi1fLW3jr4roVNFD8mU5Ah88K6qlAd5p95wQDkkr9/rLnxlT9ullmB71RsLkd
sneC3ltL2soB7caqszzdcBMq8PJpc9wZK6LApwR3OTM4DHpktLsoMfWtrrXNfx/l1zImrSrdMB9N
IPaGJtupEAK+yVdtk59wo/NAkHgEzsEGppC6p7Zx8srmJkuKYgDEHEWSqCYXm2JtjdraLi1JsHwL
BClEWb6gQNhwgI7O3FJr4fnlnqpZot4eFRushh54aUxvaINa3qHe3/wt2gecLBagY819Fyk2Xox2
ROgTIQKYgQHx1XxNaqFiUzY1AD9K9+5Hivzk2NgL8/PBaLdL0F/3yHiLr8ejbx2OBHAd7x7/lEq5
Hl45YYJNs+jsG05se6Lz/63FyAeD+IV9tWrnA109UDzY2O2sEIVUsnQoiLUKKrLUiGxnsLD7ty+W
3Cum5kN0xqRSgyp7eZpQB9Dxi3e2B/qfk1ROH9LVPZK5eA7B3wbRD6uw3/SOgQ201iedE18Wc4uU
KRJ//YuYTU0GyBbTBLQUJWJUEubP8EVQ72BUPWFtWwx3uBXw9HW5blIlAi5M6g/LjPfag6r8fhlG
GUPKDgJ+2vHrgGhEMztMIcNF2hyq2SZegr6+pAXwGusRAwvcX+WvSH8JY5z1tVaH3L5jBL+WBwOq
gB6XTUpSzK3wpkTvKTEAKwQBHU62A+gsqqjh7dNETqQCKTxj6D/SfL1qJ8qZXPFyY+JpTCBdkoRK
6B3VP3X+t6zqZU2b7M3IBPU2GUEThf0N57w7Ehpk1IUDAKn7ALndhcPkpmSQaoMi9XorCh3hPIcV
xi62fFd3zfKCvqvo6vOQTfTSwiWXDx094XGLfs8wL8/HiZbvcpy2DYKk6XRhN1dLNTG8KeYwiwDt
14NjqnnovyyuaPWQoxI4hdFvmLmr2x9Jo1LALVgKsKYCjzMb1T4+vJ10RrKTM6bYvyU0nVJVjVIF
NOydUfFqMBNzSOoS+rMCci5hjwCMtb47Bj3+S53d+TAptULnhF80gpKq1ZqqQ+nNGDejTRfUzTqd
SToIdY0WS9C0WXoEDwSBep09PDfbS+CvrlEdvM2cmDT9EHnynUP92YdbSQeU719p0UW9wcDNw/9k
NXgZc+idPZkRBc4bOn+29d+bRGY9C1NHHkCkEm6vDzIA/W2mafdgyE9/XuAk5DNYKkUvpeip2uqK
ISWkoyTnpQ+0JQz2+9iUhNBRSiawhv2mD6rhdAfmj0Qoz1Rc7cGk1LsSi4s1TUjjxluJFp8zJxfz
Ukg1/wNBR72ZFIbOY9nCSdPebbdgRP/jHgkA9P2TKuBOD3kRExK+Z8TBoHbLpowvvu9IJYGbEUFg
Pm9VFlBzFJx0QpD/rqmG6YeoOFZIG3TACdtapAyn4QmDq/9x+aZS0m9tUuuDOSanjf5Cs5AUzRfZ
oERAHBaQFsLti8VpRK/Sk/FPDHW6mGR02dq6rb8DvbcrlxodTXgSHmx3ZkU8U4nz65fV+mgmGEml
N6dnIPZhV5PDHZINSZAL6M35YXo2s4y6arpQeJVupS/ODBKAG+Sc5Ckj8QuBV0FgHBRFBlPf+oZm
/lZw5oCgRUTNtVC0IehPVn2Vxn3xkP06J/DQuktuSP2lEVCJCmyounP+IC3GlCYYZuiL6g5owg+C
6pMnMoHGZuJnL1iV0P6W3mqm4IJHfvmt6XoFl9FowVyzmOoVxMdZ/kqre9ar0kUNr3fHBp5BhPKb
09721Aebl5cJva3dMhuFuEOeGWKp+MkWJc+t7NPZJLaDNmhz7eWTgecq9YDl6lF+fs45XQRImKCY
AOabQOnqPoFReTuhR3hkI+GLucmkD3LpH2DMFo/J8Hwf0UAn9O6RbH0Tpp/Uw6BZJ/OO0CEk5PHI
MdrswJmKvgtPOcN8hFz2QK9wCKnkUvRKTzoX1l5L8NQnAZ/BQ5UxOS7ahzHodfJEMsvHN0/8JCNn
3g1v81DU9pp6SzZT2PqmmUG9sFp1xU6ro4SY+s6bc9EZfIHaX6mm7jD6EmdrY447ZX7MNEdzapK+
NbiBUiKM4nkJFy1QUlSg5umPAFpsDTVyPP1J2vnoMGJHZAyLoEHIHC3UDHqjNS8SgKkUThy+bvXq
Oa8N9dhexOLBMsMeVpbNxYr64mHUwE8fHfuT1f9KkEai6Wiq7aA5zBBdfXAFXcbBHK7ai/iK5oyw
A4HXrWXQTAAWO8zMb6JZSsvqnpAGOztAf4WbTGSsO9ymjSC+/Lv+6hns0TJKh1LiepUX7Crnexg3
Q/e/wy+IL3KvMkF0oMa0IXf+UYBplGHCNIv6pMFa3aqz2kiNFv7OFA/76Mtl1m6ustxasqkgpHQT
ktXqCGDVCYEaHzu4R+Nk+mQC/S7jIK/1ZwnF5tt+54EklAB/c+OQSNjdGNXmRRIkpjeMJLM50OMn
L3QcXIjO+zQ2aT4nGTBJPVKJxAWA1vEdmB6+QEXj+l33Yw2qE8/x9MDJ3GlUHpIw5jdgXlgKS3SI
uKU0CGnFvqSruFRuCTx+CF7oaArxyyqzw5NEgXhbAE+0viQ58eQHppQ3Z8yG2umHepcDNvGRM3oU
/LBkOrvnFWlF/nHRnUswVJDlHPALESK9TI2RNcO9FQShnx+jbIUeTod5F1/YHm8XDytGD1ZffMBY
fCfy4ngk+YZpvl2bqq4cOLlsw6EgQpEOLwCMF6IW137uxxdErxN86WnJs/2+bKQ6ylaJDvNvhWtg
IStdUKr+xJK0ThZCzmSFNZXXUjRJFu8zfXAZ4wekwV/FKU4T5l3q+EvYBkRbjWIcXxb8tmW82fgH
M/XuJQH+5aiQYIWlebNOH91ORK+qWt2PcgCmxOy6ezM/ZJlqDT8XoMnordVpf0r/0LvYZP4CCMtF
YWtQCf1/D5V0E2CAFjRf71rnK+L/qk0jmvyIX0MQZHSFL98GE1ErPSUxbnOEl3JzZonbPSZNGplB
0l6V/BowhSCrBFho7FB8bizmrrdsdlkx0SkM/9ctM5xi+ecktAbdL+Kl51tNorfIvXNzm20xAdOC
e9ADcfRtAzqDOkieDCNrYRka/vQD/T7TQcYh9KHKixT/oPfYLRWm8BMHN1iwqivut+uXOP4TLegX
BwwfjD6jFgeyq8l84S+lo+1sgzrRnvUfMp1BlDrRjXnmIlthRkxEvQVnXG4THsrXRblTcMiBX/mR
XrXiJOvuz4jN61G/XxZyeSOblfP3BE/GCRYhdntwhtRXCTh5FJEWkG9xmnqq90CXyWIMs7esfCzZ
H46HhTBb+Wc14fRDTZHaFS40iFGMG5EZEh6wV+6amY9S+5DshbctS8kvUwqm/V9cLhWihwltHgGd
9b5oktajAqZm9wdjjU40NZM5arFSOMBYV4/HqimjVRvR4EGFM67nYWXxYiNPJl+vDfbVZf3NLe6k
dGqzpVZXIRFY5nAACQQjezicrXszSbnx1rv+6eMFj+kQjuyraQMWZG2LdSb619qJB7q2T64Z+iu3
Lw34xHrmA+/KuLffPv6aGBGFZN5bBUboyr/xrrSs7OnDon9VysXEhNzPH6aWGebRB1hPNHZAIz1u
YxlVpD5lxoH3dB0xmXwjJUtX1Sbjcp/BOb+6SMClXm/EnIi0N4EtVNbi9xBfDzqH6ZTEak2UD3pQ
M/y25okSQ4+bvlZ3zXUveZhXbmKTDj3MuZcnF0yeTusrv1NSxvWxa8m1yFejhqbZfN0925SOOmH3
iVFz8/0iAvecLF2YNeMbSKU8uLmVnJpFDlsljigLugBrHKcjaxY4I6MT3DJoXUPORSEtcsAAngdl
25uRjwrIEDCow95avWb8vLwOuiXGwC/Q9fmvIgygtPR/FTdBgSdsaPBJoTj4tCMUcvQ9QcMug/Q+
7uh5Hv2uQYPznXBGAsrcQuvUT0oLWp2li/Kgghb5AlUykGWdiKZ4/oQfzpXY7Xmt/c/z5BXwOvHm
LlwWnpax65Z3KdtvYckpm/+5r4pGVzqDLJH6p7ay/mtefH9mxi2jfSh0tqNvZrkRwv9KOrXH/uK0
kpwm2VHF1yT4dK5OPC9lyghk7vtILl0vohOezozTPE1M6+ka8tf3Epi+MaovykNGWO0O6haa/SAV
IKrwriyXJUMFDCcIuRb1S7JQcL9bvm6P+KE+TfPIx4o5RHCd0YqSI3UL2DJFZYGtDX6MIWUm7kQ6
f/oCR7v7/hh7EjJK6WDkjmWrKEVgn5EglYUTk+O5Zq/M8I+ZWwfSLII3vCt9J91gGogvMMZI8JI7
wauJYbFCMn5RIml2PPZ0oCFJGd58oWCODiDd7IyxoZuWeVc1uMQUiQgIfzjXvjI2ILgfLu5FvSt3
Z5phPy6xzJwjaG3deQI8NU/XjwXJ3Dc/3ixvCKYrZIxvNf7brGUC6UuIJbgabrftqLddDT46jToZ
/i67EX6qXXI7zdCs52XIk3xyK4WZQ7t950eS72EcNgGQGDWag1kEpOWnnGpJvNayiO6yupIb54WU
fifluvsC30bjDAy6txyjFmab45SPy97qskIH82fBWIwKWnExgR/rq2cTaDi/4lD85T1V5gUwFt+z
3LanwjY8C2etJ/H4qae/4UCdMYJtGLROavwZk6Hrwu4ccdaN984JABUjBVhNsEvg9OzjhvCB6pf+
Pqtsa2Z+pyu8QCckSpuoYL9li2NHiCqqod4IG8s23FeDYMgSoOLnoHE+PPwnIn98TgOxiKNG9nCi
kCU0Nf1FzpMMk2I2YwAhTVyWRU95EQ37bVoleSrXterJKBwwDqfkRcoMuzwUAvSoLaCwJSBLGcI5
3m0tC5/aVamPb0imtI/vLQcXQMenTWhHWAWX26STKTEEiBFZzLYtyq6oMa6j95R+bZZwn/ZprCVw
r0NHQj/x3K/Gq56Mg4ecGPgXqcAm9Z6FRBd8CFhjXKO2FuGPuCF43OV4fShY0U2DR8PYQT0mo+sF
t716bBbMOym+4VMj12usZx4PCYqJWEa9mEGU2RbiwkbJZ/KSLW3Y/JjqEHuG2vstBl1ypiS9D47F
pfbZ9a6Vnh9lWpvZ4qxm5DHfMfWLZRl16JfxT1IShXKG6bdfHOBazcZxtLT02CAxKtxs/YgFVYLb
uzmevDJcCZP5vl8YvXbaZPhWpSEzEW/RZ2kMbtSXaseVRwtTUGWWpptH9L58bApeCpds5z5B80OE
6fp1ZRuR2IAzDSL5lKrXVxbse3moHrf/GNe5aUDmKpucv9xt7jdPGtTTnocHFutq0muKJ3Lq/EM/
av04+Q3Ttf3uHmW6+2Dt24/hvHYwFQvQ8EB1v4B+zkyZUbkRlVk4bGAg8DOuw1oBS/McqJaU3D/q
AVr8hUo3EX2vpf3DQxFoHsa8Nr6qKQK4AzYYe+oK0dNs1484XDJObdwmyYzYE95GTeDS5lCd+4s1
z0exm0p82kfdbxzwOg8SvO3LN8RjM32E9V6X8+fy9MlVJ0otAAv4VnKYKwE+IrX4ZwBFPamg7tME
sewyJS98XCVDXN1H0/dVH71ewwTKDTaNU92NSlRNfDxrwuoRyfYwpG/LC/6Qdlppwhd+Pe0xNy7j
tpSn5XhPZVfDHTGyUc19C7jmhOdKWg/BQQFINgencoOOTvW4jmOoueOGtmDhjJkBTswW9R/iXFox
IzhRCvcGmIAUyMpw+sL2a+sY+IkUi2Kq2r6j33G+j4D+Qya0ucXZFldMPh4lBLba9kGyGU+zQIEI
kbQ9YCA3WOI1LcQuTj8WPE+hO1r7OgIunoANbsJqnNV5JtWJ2u2OJ+466tRU/cUtbI1vHCaBUiBB
EjLMmhNeot9p9+xzL3l/nW1x3PQ1Dy5eaw/L9MWe4z4bKZxHCiKgadsksj7RS9zzhi99u+EN4Omc
R4NPweSX8VhOkS4j1j0rImmEjaSXOt2q/OQ5uHSIhZxf0hfJqeNRw21nvY+RK22AzIpNPPFNfOoO
zKnDUbyjzUHEIkXz1UPPWmEeA3GjDwyesp/s22C497/rOFm5notUHGNJLdA0Rhvn7DnA++v0rUN9
s1XRm1kew3kOgj1Qn21tw4fCOXkhP7B30qf9UK51bFBVlb8ziNKpB9fxodyxr7wCwS9Xg4WpLpZL
gKw2F2t8wVSeVJFGj5UqKVJVZ7OTC+LLqDJ5MhrSGS1p2B16k+KKoJmk9FUFIKWwGJ2laED+hk5w
m+u/TJQwVZVchfVoCz0qkKl26NcqLclTK6FdzRw4aGJd8V7ktp9+TyPgiKIkwspuqoK0CE8jXTH9
NfHmK19STrdGFgT/Y6XsLoo72eKzrQRFsqu5DGi3RZ/CGEz7q//E0celJqh7WOiLmwyyLqEOApDG
zpLKFY7Nw0BBG15HX9AATonKZElb4IE9pqOEnJf68juA7VnjCJeSdH3i2HdiyFFdr68tFY2HzhmR
Tvxv7MEAyGhLxfnWFAFsZjCL19tMtEp7c5qV0MW7Pw7sEWACm5zoQU8Wc3bDgiQxiTNZcWm3PF90
LEPUNcq1lJPY/fmKHFK0NHpBwhuVZrdadoOq0oUAY/BTvXacAieeqixXZ9tDGUyOkh77pIHLamRS
QUgGvaKRucY7L/rvSQuTm9FJs35eyNvFVs9ulBQURPxwEz9cPDnerO5Z38hcgT3xwOzQLa8huuZL
MoVrrZkLb3mT9ar2LdcTpD9ODw+GyhFcNcFdthPgE2zZLmDLkWN60ozCLuEtrgfHUvcqHoQmGV7L
NAlKKxqFcBIZcK1RqrekD/pd1DsO52cGSrG1JZV0KsG88praSJAdXVeJJFxqLjLLpzJPs7lPNyau
fSqei9FKjZCgU75J6RDebzioOFQrt7XAXZyNQmK+b6CtgED917QQJLYvuj98qv5bNb2LHJKd2IPE
4elCm+bQni+ggq2GHs7QYrh1eVFigUSZGJtmngsM6NhO+JVTPecm4Sc1BI7WuOaLPHQ2tZXIoKom
6a5QRA4sKf6fHd/6T+O0q+4RFl2VJhgCCrcWDVLsKVYhcP9NQWwZwRrgoCLIXHmx2vKBB3tXe4XF
TMrDXG3d17Sx43ouO9eO4uaM1RheDztyyTp0uoYmS1JFs22g/DWWHotWSy2TI656eSltf2JRHktY
Sa5YpPsSeE7+omLQdr+t5LVxhBAMIQnDgpG/GKEhFJbYlJlGBq0h50Qn3aIFYO45PyWw2xpUC7/v
TZzu4vpKoBwErYnJkR9aZI2tUosyo2VG3blOikPfUV11TwnZQ8OLi6W3Qr/g8i4n0ueO4rEfDAOL
iIlircIQk+ZRITPgtGgZOGLqpil1ss+ISm4h6SsgDgbhorAs6OuGwl4m1IXjJI7S9sm1Ej2U/nCm
7idAAPBSPiw6OXCuqlG8DqhBwhYm+IUKOISucCQuYM9ncMEtCOOmh7Ww6fzfGxrKmGo3B0wwshSE
tH23evLKJnXOhfMwwFMsnWMMUUpTj991LZaWl7o4eSRAjoVxGl13wUjSiQOTUtO22MMJroe8Xc2Z
yItu13vnnhTcsOUa1OMbC0TxBtUZ3Ihk/7j2F97Xyq/kBHbME3afa5azkXkPNOgH9JG7C8LLwgOu
S8xeLFA3SiUJCjjVclPTdi7zHFukDmoEfoE5MzVDdE6ijUwF90KlkoZzh8Q0nL1mya+7pC6TvoTy
OnVw494yoeoUmNZ+OwspXniCeWzLu1C/8IVqtgTt5d3YzPrI+u82Rn7RUuiFdliXfoy+wPPbKVje
IOGgAvI5S0o3je2uE1Hnt2/OGdBGtTRYN2L73XzHEQx3HX7jaKfivWJtSycU6bDx6zWd+iSCwOpP
LZcyr0mC5PLS/3hsnfSBMs26TN8Zafw1TKl0nhwdZAyWjhofoKqtNrNXxszIhGgCH0QiIwbjNcVX
ExxcRKsfRyHkwgAk7QalyaTl75lIB2vO+IV6JBKh+8cz0Olzlx/Flc7dSoZo8Gah1i9aeAoE+wS3
eCqnpGLT2DADxGM81jKkKBR+Lqvh0Yht1rHBger9w2Ke2/2abKPuOL90fCDoa/Di/cYV4ld6JCpS
aPAIhbFzWzGT90kqip1X4cy4Xau2/CzQXRFtaxHXt4Iz7eGy35OG3NpKmMkBfKoNpO8tVIhkhZS+
a6YmVtEbHUCNIKCCDuUf3dNcnCQ0zkeZguwR6OT/I+33lYV7HwmqkzNhh5kRNOgsNSHiQX1bS18g
TFF6l9DAobsD9QBOq/FDzclLzfJd3MwpLsDInE0viLU5O6+ydrBb/KgPpJ78xxbYFv2z+P0OeX9j
4FuwxtWPtMnr4A741o4eMxBX+kx1j3pgxBEe1tOrVTBtdJS/iDE0Gv1hU0TnJMRoPqcsZif4M97o
7SZ5a6FRjx9mGP53yzLC8JbAc46h5jjRvZiyqnlCpED9cP6cUGIXwmRkLspog1jXRvSCEr99tCa8
JzQtgOZu/uA9n+KtWTTtouMqBXZt3NsuDHgzzFefBAss22LZdy+YDaRRK8HI2oVWoKhQt/GNE0yu
sJ//u0BzLLCrnfJLnJ2Y2ZMh+MDqYYPMALcGyXvueZi6F6osRPrfL1BmScXpajxq0v4Yrxk6pM9w
wo1XG25wjs3bNOUufbWfIrY+Ce+dcpUVcWbDLIWznyglKbYfhekjJe/KsSP5J8zEhpwYOs5HQ48e
kUgXo3m/rgABbcwjX/DikKKKCSR/1JDQdVybydV/lBgnDNsx+ZWSWCjKYBGG8ouGeLvg+S7//xW3
A9Z5i0QBcN/YnFPqLjLYrSZbyBgp9OvxPDWaBg6RXqW2S8zafo41FzaxWghBIPrjHRju9KYXJ2ah
gcRqjOWER7s+sDOdGYAx2IDuUpCyu82nzdOAlT2vx5o9YqZLyDZu4FMaKOFLcOmVroV6MKm4zGQM
0VCPHffYJAFtFZzRhCLxKUa43ZYfnH5XghS3Yoyq7N+90TrwvKvhQJLHFUs2gRRBF0Qrgb+sVK1R
17VXnir66SjEdoWwhswrdU7OW6DHKQVrMbzotFhXNgUGKezH8k0jL/c60uQhT4na7iBFEHdDFyIo
C8vGkjF16Xb4eZLxvQ6UqJo32i1zlffsq3Z4bHuCbbcMA1z4em7uiUyrH0D/MJtuWFptRyzDtV6x
lCzK7lsNtrvLzcQ4n7WWM5WDWEtrhYPACNT3bMx91ciaH4kG96Xu8hgwvozWJZDVb3H2JvHqd5ND
fDbTm/cnqc2CU6tX4nE0z7xS87tAzA2yISM3FmfXmTjU+VDNouWAmGxdpkJYjP5XpU95z5jr6KDu
iCgjRK1sQEe1OxZ4jTyjLiE/cJvk9XM6mjlG3RCb9CLQ5drX67GClXKZAcsyRwP04jasogPI7+dr
SKguYucmsDnyBGdnEqNVCnLdq2zrV7Ftu5uqd46t4b4gR9sl53/qN9FyrILPg+VCicNeK+gEuJWn
2OgiKOm+vfnwusInxDTEMcX5Qa1MQ4d6FrOdNC3FBbjDvAsA9IOExogblqVfxjHzz3BFfVuQjUTo
Hwhw4zDDlY7Z9B5yoSKn3seVwqy7ukw7wiG+T3uyrdlHWtDLBNmzQHSDybw122YUzCy7qU5IBUSW
uN+LrznWN4W3PCvNgFR/zxKPjK503SyOEITV20ZdsJQuZLbjw4xpmAEGlJ6n8bjC5r5Yrh1ac+OV
LY8Y6fJDCjazATJidcOWli+DUgycrFGlT714x2vKU2W7lIre3gUjEf9MV9FnGMZc+Ad0x3IF8o1V
Ur1DFYsYLs0CCf7ZADia1cHjYaQGYFawoTdIfbWbEZajRpkQZx59anCRBIGzroZ4gW5Wht2CATq/
n0G0yUiPma0GK5r6t4pfSYvg0oHWyJ/VovOJw5lzfLv6Sh5ih3/Qna4ek/DFu2OzOBqTnng3XlMH
Z5VWoyWyG/JyW8aeByhdBOi0fWPMI0rI/S+c1mHPS1vmOZvNBphUf3mDbe4IUWhFvEZfD6P/+J78
eMf+erACBMlgEZBkAx2sYzPdvHh2PSI70fU2JOzkNWZivLDx3qWmL8vRAUXGI7BS7t+yXPnaeb+V
0e3/NEJnCDKYzG/PX2TejsjeG1RGh8qqEhQMxHD4ttjC00In0Vm3Fl6TZNQPpXCQsv12/t2/b3Yl
h5RYaCC11YTUtjXKgunZmo8fbkl24KmtU5D6zo2X0vsFG+tNLcwgHo5JSTUiPTUZsH5UA7H/KQLs
o2OI0q9XnsMnaI5MZOq4tbpFxOjqcdKajbU4QhrrbtHaZDtF0nqOosRgXYzcRx4JgKiGy4uM1PqA
51UodS7M1HBPrA/6l8ST71jp1E4mTQnaEYiYVTGPXmHzawn6gUnCzQ2WAk+mTHxY2QH3r54jZChP
LB8LAWOckiWJXx3ICdC5pR8QRhj9NjLqpYigL1GWDKk0E0wgv7Jd/ig7S7v/EAjcijHvKgFj+Zzq
Vi5yM7Knh/XTHUdljRw6AQ==
`pragma protect end_protected
module DVI_TX_Top (
  I_rst_n,
  I_rgb_clk,
  I_rgb_vs,
  I_rgb_hs,
  I_rgb_de,
  I_rgb_r,
  I_rgb_g,
  I_rgb_b,
  O_tmds_clk_p,
  O_tmds_clk_n,
  O_tmds_data_p,
  O_tmds_data_n
)
;
input I_rst_n;
input I_rgb_clk;
input I_rgb_vs;
input I_rgb_hs;
input I_rgb_de;
input [7:0] I_rgb_r;
input [7:0] I_rgb_g;
input [7:0] I_rgb_b;
output O_tmds_clk_p;
output O_tmds_clk_n;
output [2:0] O_tmds_data_p;
output [2:0] O_tmds_data_n;
wire VCC;
wire GND;
  \~rgb2dvi.DVI_TX_Top  rgb2dvi_inst (
    .I_rgb_clk(I_rgb_clk),
    .I_rst_n(I_rst_n),
    .I_rgb_de(I_rgb_de),
    .I_rgb_vs(I_rgb_vs),
    .I_rgb_hs(I_rgb_hs),
    .I_rgb_r(I_rgb_r[7:0]),
    .I_rgb_g(I_rgb_g[7:0]),
    .I_rgb_b(I_rgb_b[7:0]),
    .O_tmds_clk_p(O_tmds_clk_p),
    .O_tmds_clk_n(O_tmds_clk_n),
    .O_tmds_data_p(O_tmds_data_p[2:0]),
    .O_tmds_data_n(O_tmds_data_n[2:0])
);
  VCC VCC_cZ (
    .V(VCC)
);
  GND GND_cZ (
    .G(GND)
);
  GSR GSR (
    .GSRI(VCC) 
);
endmodule /* DVI_TX_Top */
